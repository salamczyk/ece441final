library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package project_package is
	type weight_1 is array (0 to 783, 0 to 127) of integer;   
	type weight_2 is array (0 to 127, 0 to 9) of integer;	
	
	type intermediate_output is array (0 to 127) of integer;
	type final_output is array (0 to 9) of integer;	  
	
	type image is array(0 to 783) of integer; 
	
	constant weights_1 : weight_1 := ((17,6,-12,-7,-18,0,0,-5,3,-15,9,-4,6,-19,-16,-10,-16,-20,9,-17,1,3,18,17,-13,0,-4,1,13,9,-11,-13,2,4,4,-4,-12,-2,-13,-16,4,7,19,9,-16,-6,-3,14,-5,-9,-18,12,-17,0,-2,14,0,9,4,14,0,-16,-1,7,5,-10,11,-19,-15,-18,-15,-10,6,6,19,-12,6,8,-16,10,5,15,2,17,-1,17,9,-20,-7,8,-18,-14,-18,1,15,-12,16,-5,0,-8,15,11,-16,-3,-5,-12,-12,-18,-19,7,14,-2,8,6,13,7,7,18,0,11,-10,0,18,-6,17,-10,-13,-19),
	(-19,-13,-15,-17,0,11,4,-8,-17,-14,-6,-4,11,13,1,1,-7,11,11,-5,7,11,4,-13,-9,-9,4,-3,8,-6,4,-20,-12,-5,5,-9,10,-3,8,-14,2,7,14,5,3,-16,-15,-12,0,-19,14,-13,-15,-14,-18,-8,-13,-18,-19,19,-7,13,19,-8,-15,1,-18,15,-16,0,2,7,-5,4,-7,-1,15,11,2,10,3,-1,1,-4,-9,-14,-5,-6,7,-9,13,-19,-19,-17,18,-14,-3,0,-19,8,-11,6,-5,-12,-14,11,-4,19,-2,-5,12,5,14,3,4,0,19,8,-16,1,1,-7,17,17,14,-5,5,0),
	(-11,8,19,-5,20,18,16,-17,14,-19,-9,18,-2,-1,-11,17,10,-10,-6,0,-20,-3,-5,-9,8,14,-19,-17,-13,-2,-13,0,-10,17,-13,12,7,-19,-17,-4,15,20,8,-12,0,12,-18,17,3,2,16,6,-8,12,16,14,-19,-11,19,2,2,-2,16,-17,9,1,-8,-17,5,-5,3,-12,19,16,-6,13,-4,14,-9,0,-16,4,-4,-15,-20,12,11,0,-5,-13,16,-3,-17,6,-14,16,9,12,-11,-20,-2,-15,-7,16,-17,9,2,2,-6,9,0,-14,-1,-7,17,11,-17,-7,12,-8,-1,14,13,17,6,10,16,-10),
	(6,-1,4,-16,-8,1,4,1,-6,13,15,-14,-15,19,19,-7,-12,3,8,0,6,-10,-15,-20,-19,-2,15,15,-4,-11,-19,20,3,-19,-15,-1,9,15,-5,-14,-9,10,-9,14,14,2,-16,4,-6,10,8,8,16,-12,-2,-2,2,-12,5,-19,1,15,-10,17,-14,-4,18,-8,-13,-18,17,5,-2,-2,-3,-6,9,-2,-16,-14,-3,-4,-5,-16,-1,-14,3,-5,-13,-1,-16,-2,-5,4,9,-16,-4,0,13,10,18,7,0,-3,10,0,0,-8,-8,18,9,-9,6,19,19,18,-5,-11,0,-15,11,5,-9,-3,2,5,-8,-15),
	(13,6,-9,-11,8,1,5,-9,0,14,-20,-15,13,6,4,-2,15,0,11,-9,-19,16,0,-9,-16,17,12,-2,16,-4,-2,9,-4,3,-16,-16,-10,11,13,8,-15,17,-2,-4,-13,8,3,17,-9,-4,9,-9,-9,8,12,1,0,19,15,17,16,-7,16,3,-20,-15,5,10,-10,-12,10,10,-5,-6,-12,13,-15,13,-5,19,2,-13,8,11,18,-5,-20,-10,15,-3,-1,-10,3,11,-20,18,-16,-18,10,17,8,-18,19,-8,14,7,14,-2,20,5,14,0,-5,-2,11,19,9,-15,-17,-4,-5,9,3,-13,10,0,-18,4),
	(-13,7,-14,-7,-3,1,6,-1,-19,-20,-3,-18,20,2,10,18,9,19,0,17,-11,-1,8,-11,2,-1,10,-16,-13,14,16,9,3,10,-7,-15,-1,-9,13,5,14,5,-16,-7,-13,-6,15,-11,-3,-10,-15,5,-9,-2,0,13,17,-20,7,13,-19,16,-9,-20,-6,4,-17,3,16,0,2,-18,-6,1,-18,-13,-14,7,-14,-6,3,-7,-12,-10,19,-17,-16,12,-15,-5,4,-12,4,12,-5,-9,7,-15,-2,-5,-19,-11,-10,-9,-7,7,0,1,-17,1,-1,-4,20,-5,8,10,-3,-3,-17,-8,-9,-13,-12,0,-14,6,4,-17),
	(-1,-1,-3,9,0,6,-15,0,1,-17,-11,11,3,10,3,-19,11,9,-18,10,-2,-12,17,-18,5,10,6,-8,-3,-5,-10,10,-10,-19,-20,7,-6,-8,0,-13,-14,16,4,7,12,-5,-14,19,-12,5,-15,1,3,-8,16,-16,-11,13,15,-9,7,14,17,0,-15,8,-9,-7,-16,-10,4,-3,-11,-6,-8,-2,-18,-13,11,13,-14,-11,7,9,4,-9,3,-12,-3,-16,15,2,-11,-10,7,13,-5,-5,5,14,5,-15,-10,17,-14,14,4,4,17,-19,0,10,2,0,5,-1,-18,-15,-18,-8,14,0,5,3,-8,-4,7,5),
	(-8,-16,4,10,-13,-18,19,-14,17,-11,-9,2,-3,-4,-5,10,-4,-9,13,17,17,-14,-4,2,0,-11,5,-4,-10,-6,16,-9,4,6,-8,13,-15,-4,20,15,-15,11,-12,-16,1,6,8,4,-9,-2,-8,-7,5,11,11,3,-19,0,8,-12,16,-15,-20,-5,14,10,4,20,7,-2,-2,16,18,-8,12,-15,-19,12,9,8,12,16,-11,-11,-11,-4,10,-2,-18,-4,-5,-7,-19,0,9,11,-2,-17,-2,0,20,-9,19,-10,-20,-11,-4,-12,-11,-12,-17,20,1,-13,7,-7,13,-1,5,6,-19,-5,6,16,8,-14,3,0),
	(-14,-5,11,20,10,8,-14,-18,9,12,-15,13,11,3,0,19,-20,-17,7,1,-20,12,4,-6,8,-19,1,-1,3,18,14,2,-19,2,-4,-5,2,1,20,15,4,-5,-17,10,-19,9,-16,-8,-12,-11,19,20,-18,1,11,12,14,-4,17,-2,-8,-13,-4,-10,-15,-15,-9,-14,1,-9,16,-4,14,-20,0,15,-18,-16,14,0,9,-4,-16,-20,6,-11,-15,-6,15,-11,0,11,-19,-11,-18,-7,2,6,17,-8,0,-5,18,10,4,-15,-10,8,8,20,-2,13,-16,-19,15,10,-12,-8,14,14,-12,-3,-1,4,-4,11,-14,-7),
	(14,-1,-8,16,-2,1,15,6,0,13,11,1,0,-17,6,13,17,16,11,14,10,-20,-2,9,-17,4,-4,-2,-4,-9,-4,-13,0,16,-14,15,20,8,-6,-2,17,16,2,1,1,16,-8,-18,3,17,15,-9,12,19,-9,-9,-7,5,-10,-18,-16,6,-16,-7,20,12,-18,19,-20,0,1,5,-15,-18,8,-15,-12,-16,-20,5,11,-17,7,3,6,-14,17,7,-2,9,-6,-17,5,-17,4,12,-20,8,10,8,17,18,-3,-19,10,-11,-4,10,2,-6,-8,14,-19,3,14,6,-5,4,-7,19,19,-4,4,6,-14,-12,-16,-1),
	(-16,0,0,15,-1,6,1,-11,-5,20,-9,12,16,-10,-3,-19,-10,2,13,0,12,-9,9,6,10,2,19,-1,-10,20,12,-15,-13,-15,18,-11,-12,0,5,19,-1,-6,-18,14,-3,-4,16,-10,14,-5,12,-8,5,-5,-17,14,4,-12,16,8,-9,11,14,20,-6,18,13,4,12,10,14,0,18,-5,13,-10,10,0,-14,-18,15,-6,1,7,-17,0,17,-2,-12,-18,1,14,20,3,-8,-1,-3,2,-16,-7,-14,4,8,-5,-10,-4,-15,15,-9,11,-3,-11,-20,3,-10,-13,0,-4,-20,-6,-17,-13,17,-7,8,-3,-17,-9),
	(-14,8,-18,-12,-16,-14,-18,8,-20,-7,-12,6,-17,17,-17,-13,9,-6,10,11,4,-17,5,-11,-5,-14,-7,20,9,0,17,2,-1,17,-16,11,-5,2,6,-11,-4,10,11,2,-3,-8,-7,-12,0,-3,0,14,-16,8,-6,-5,4,-18,-6,-2,-3,-10,11,3,-12,16,-16,12,16,0,11,0,19,-10,-1,-12,3,0,18,3,-12,-11,19,5,15,14,14,11,19,8,9,-4,0,7,8,14,1,13,11,13,0,15,4,3,6,9,-8,12,-12,2,-20,9,-19,17,2,0,8,1,13,-7,-18,-19,-4,10,0,0,-13,-7),
	(7,17,8,-12,11,15,9,-4,6,15,-8,28,-2,13,5,1,11,-2,-17,-15,-16,-18,5,-1,7,2,8,8,-6,1,-16,21,0,34,0,-8,16,1,1,-7,14,32,-6,8,-24,5,-1,-3,-20,13,-5,5,25,-12,6,-17,-1,2,-15,6,-12,9,-6,12,1,25,-11,12,-3,-5,-12,22,-16,0,4,-10,2,1,-5,-18,-14,-9,-33,15,-24,19,-18,26,-6,10,-3,1,19,20,6,16,-1,0,0,-11,20,13,-4,-22,-11,-7,12,22,-9,-24,2,4,-2,4,15,22,18,-5,-8,-18,-7,7,25,11,-13,-5,-8,-14),
	(14,12,-21,-6,0,9,16,-20,0,6,8,17,10,-7,11,-3,-16,-10,-1,6,17,-1,-13,-18,11,1,0,26,-6,0,2,0,8,-3,-9,12,14,-16,-19,-13,8,17,-8,3,-13,17,-4,13,9,20,-6,8,-9,-32,4,12,0,7,3,0,20,4,1,-18,-4,0,16,-4,-26,9,21,1,1,-16,4,9,-20,25,-21,-1,-7,-26,-7,-2,-10,-17,2,14,29,-5,29,-3,9,-3,-8,-12,-2,-5,-11,2,-2,31,3,-20,-12,-14,-13,16,-4,-23,-7,-1,9,5,6,18,22,-4,17,-2,14,5,16,-19,7,8,8,-9),
	(-8,-35,-2,8,3,14,26,-6,13,-16,13,-5,-9,-6,12,0,-9,4,3,0,-8,5,-17,0,-8,16,17,2,-19,-15,-6,5,-4,14,10,-16,21,-14,-12,11,-16,-23,19,24,-6,-18,-2,18,-14,-21,4,-8,15,15,20,7,-20,4,-23,20,-7,1,7,4,7,-20,-10,-9,7,-12,22,21,2,9,2,-3,4,15,-22,-5,7,-5,6,5,14,-4,19,6,10,19,8,-10,-5,28,-8,6,6,28,-26,1,3,11,6,-5,20,15,0,9,14,-15,-14,-4,-13,6,16,32,16,20,-12,-4,20,-15,23,11,1,-23,-9,-13),
	(-12,6,-18,18,-23,8,18,-13,-13,13,-2,11,-9,-13,-20,-10,1,3,-14,-14,4,0,-24,-1,6,13,18,20,19,-2,0,-18,-3,-12,0,-5,13,13,8,13,8,16,10,20,13,-1,1,17,0,14,9,-7,-1,2,4,-7,8,7,-6,4,-8,-12,15,-18,12,-15,15,9,16,-19,2,-17,-8,-18,-19,15,18,7,0,16,-16,2,-15,-23,6,1,10,1,-6,-18,-10,-1,-19,-2,14,-5,-9,14,-20,19,11,-7,0,1,-13,-16,-2,11,12,-12,-6,5,7,-13,4,14,4,18,0,2,-9,8,-8,-11,-2,-6,6,9),
	(-10,5,-10,14,18,1,-6,-6,4,15,-15,-20,0,-13,12,10,6,13,-15,-8,9,4,-18,15,-1,-1,5,-2,20,-5,5,8,-14,-5,-1,-10,2,5,12,-10,-12,11,-18,-2,-6,1,19,8,5,5,-6,-1,16,20,-6,19,3,7,3,10,-9,6,-2,-19,-9,11,13,-17,1,-3,10,-5,0,14,9,-3,-5,2,-14,-17,-13,2,6,-17,18,-11,-10,9,0,16,16,-12,5,14,-9,10,16,15,8,4,-5,7,-11,-4,18,18,0,3,6,0,-18,-11,-19,18,-11,-4,-19,-19,-6,-3,3,7,1,16,-14,19,10,10),
	(5,10,1,15,-2,-1,-6,-20,3,-2,-10,0,4,-15,-4,15,-8,-17,3,18,-6,-8,-7,-14,-5,2,0,-13,-3,10,-6,13,-15,8,13,-6,1,8,18,-6,0,-10,-17,-1,7,8,13,-7,3,-8,-18,9,-18,18,-6,17,4,-19,4,4,14,-3,4,-17,0,0,4,4,-15,6,-15,-3,2,-8,-2,-16,16,7,-7,3,-16,14,11,-14,3,20,13,7,7,4,-19,-8,4,10,-16,6,-20,-20,16,-4,-15,12,-20,5,-18,15,0,5,-2,14,12,-19,3,20,18,-4,0,-17,7,4,-5,-19,-12,-17,0,-16,3,-15),
	(7,-19,-1,0,7,4,10,14,-9,0,-2,16,10,10,-2,14,-15,5,6,13,-13,-2,-13,8,9,15,16,3,-10,0,-20,-6,12,2,19,-7,-15,-8,18,9,15,-3,-13,-7,9,2,7,8,-15,9,-1,16,-11,20,20,-5,-3,5,-9,8,-20,12,6,-6,-8,-18,5,-8,-5,11,-4,8,2,-7,-8,-18,0,-8,-14,-10,-6,12,-11,2,-19,5,6,-19,-6,-15,-7,-9,7,-13,17,8,19,-7,-13,13,10,-1,-13,-11,-15,-10,13,2,-1,-15,10,10,-2,-10,-5,2,0,1,-20,-19,1,5,-11,12,-12,4,10,18),
	(-6,1,2,0,4,5,4,1,5,-13,3,2,-16,4,13,20,12,-19,18,-19,-11,-10,-18,-20,10,3,-4,-9,9,-12,-5,-19,7,0,-12,14,3,19,0,7,-6,-9,-10,-18,8,4,10,10,11,5,15,17,-12,-1,11,-10,-7,-9,16,-11,-12,-18,0,18,-6,3,3,-19,-2,-4,15,-10,13,13,15,2,2,-11,-11,11,8,-3,-3,13,-10,-12,-5,18,6,10,-9,-19,18,-16,-1,0,16,19,6,20,12,10,-12,6,-2,5,-9,17,3,-5,0,-9,-5,0,13,11,-8,8,12,11,-10,8,17,20,-14,0,-8,-5),
	(-13,-9,6,-10,-3,-12,-4,-10,-19,-17,8,20,1,14,10,4,-7,-11,2,17,20,-3,-3,13,-1,-8,20,-1,-9,2,8,4,12,-19,-16,1,18,-3,-16,1,11,-15,14,2,-12,6,11,-14,2,0,-19,-18,-4,12,-18,10,6,-10,15,0,10,0,-15,3,-9,17,15,-11,-17,-17,-9,9,-5,5,14,-18,-14,-5,16,-9,-2,10,-6,-9,-6,19,13,-14,0,-9,7,-5,-14,-12,17,19,11,6,-6,-19,-11,8,1,-16,0,17,0,15,5,-12,-6,13,11,-16,-6,19,9,-2,5,9,-9,9,1,11,-14,11,-15,9),
	(-1,-5,-2,4,-3,7,-3,-18,10,-14,1,9,12,-14,20,-4,14,13,-13,17,-2,-9,-8,1,-19,-13,-17,-19,-3,17,-6,7,14,5,-11,12,0,-8,16,0,11,-12,12,0,9,-16,-13,5,17,8,-18,8,-18,-9,20,-1,-12,18,-13,-7,0,-16,-20,4,7,6,5,6,15,10,-10,10,-17,-1,-19,-7,20,16,5,20,-17,13,2,-18,-6,-3,-7,4,-14,-20,11,-2,-4,-11,17,-1,-17,16,16,13,-1,-8,-10,20,-18,-10,15,-13,18,-7,4,1,-1,-9,17,-2,9,-4,-14,-18,0,13,7,12,-17,20,-2,0),
	(-2,-7,-5,1,-14,16,-10,-10,-5,-10,3,5,-17,12,9,-15,-8,0,3,-15,-12,-17,2,-5,0,-12,10,-8,4,-7,0,9,-1,17,10,-9,0,-10,5,2,-3,-11,-5,11,-7,1,5,1,-2,-19,18,-3,-8,19,5,3,4,-16,-5,11,-17,8,0,10,-2,9,-7,-19,-20,2,-15,-6,1,-1,-3,1,16,-18,12,8,2,-5,-12,-20,2,20,10,5,-2,-5,15,-13,-11,-10,18,-13,-11,-8,-9,1,3,5,-15,6,-10,11,6,13,-2,2,-4,12,-11,11,5,-16,13,5,0,8,1,-19,-18,8,14,13,8,20),
	(0,16,-14,9,4,-3,-12,12,-4,-1,-15,-1,-14,-6,16,-7,8,9,-16,-9,-2,16,-4,14,7,13,-2,8,19,13,2,17,12,17,-3,-10,-15,6,11,5,20,20,-7,0,-14,2,-4,1,0,4,10,2,-15,5,-20,14,-11,-13,-9,-9,6,-14,8,-18,17,-16,-11,2,14,-9,-13,5,-7,16,-6,6,9,12,6,2,-5,7,1,-9,5,-15,-8,11,15,-12,-8,-3,3,-9,19,15,9,15,0,15,-2,2,-12,9,15,19,16,13,12,16,7,16,16,-20,-4,-5,1,-15,-8,0,18,6,-10,-3,13,19,-1,20),
	(-8,19,-3,12,17,-3,14,1,-3,0,-20,-1,-18,0,16,-10,-8,-3,-1,4,-13,-15,17,-1,-14,5,-14,18,15,-4,14,17,-4,-15,17,9,7,-19,-15,6,-3,-18,7,-12,8,-12,11,2,-17,6,-7,-13,-11,-12,13,15,-9,6,1,-3,8,10,15,-15,0,3,-11,20,13,-9,17,4,15,-9,-9,-19,-5,8,0,-11,12,2,-12,10,7,19,10,-12,4,-17,14,20,13,-20,0,4,-2,-9,-9,0,-5,0,16,-12,-19,2,-17,-8,5,-11,-19,-8,2,-20,11,7,-12,-10,-3,-18,-13,0,0,5,-11,13,-16,2),
	(14,16,15,-13,10,-15,-8,0,7,-14,4,17,0,11,9,-6,-20,-3,1,20,0,8,-4,-14,-3,-13,-2,-5,-6,0,10,14,1,-10,-2,-7,-13,17,-10,10,2,17,0,19,19,-7,13,4,-7,2,17,2,-2,-15,8,5,-13,13,7,-11,-2,-8,0,-3,-12,12,-19,-7,-5,5,-10,9,9,0,2,18,5,-12,-3,-20,-16,-13,2,-6,-3,-20,-20,-5,-7,3,-18,-12,10,16,13,15,-19,0,15,17,6,10,1,-11,-9,17,14,-18,16,-8,7,15,15,11,1,1,-14,-2,-8,3,-2,-7,-14,6,15,-13,-13,0),
	(12,-4,14,15,13,-6,-14,-13,-14,0,7,-3,13,19,-19,14,-20,1,19,1,-3,-1,-10,-6,-7,17,-7,10,-9,-17,7,-18,-9,-3,-6,19,16,-18,13,-12,0,13,4,-10,-11,-10,-14,8,1,-16,-11,-18,-12,-19,8,-17,4,11,16,-13,10,19,-17,0,-20,14,7,10,-13,-16,-5,13,-10,3,-9,-16,-12,-14,9,2,11,-17,7,-16,-19,16,-7,15,0,9,-16,12,13,6,13,-8,-8,-2,-9,-7,11,10,8,17,5,5,7,20,6,16,1,-9,-7,-13,12,-18,11,-16,-8,8,4,0,20,-2,7,1,-5,-16),
	(-14,-10,20,11,-11,8,1,-17,0,4,16,5,-2,9,1,-12,0,3,4,15,-14,-4,-5,19,-19,4,-15,-19,6,-4,-19,-2,7,-7,4,15,19,-14,20,15,-20,6,13,7,0,-12,5,18,-7,-17,-10,17,0,14,6,18,-19,18,20,-14,15,19,-9,14,20,-10,18,9,9,0,-6,20,11,12,-14,-5,15,-9,-20,-4,2,19,13,12,-15,-20,-11,-8,14,-1,13,11,14,9,-19,-6,-20,-2,-5,-18,-10,-10,0,-11,-6,16,17,-2,16,-15,-17,20,-16,-4,-9,3,-13,-11,-7,-6,9,5,6,-7,0,-5,14,18),
	(0,3,4,4,10,15,14,9,-12,18,11,-14,-5,-15,0,-7,4,11,18,6,-4,-1,-7,-11,-8,0,6,-13,1,-2,7,19,7,13,-1,0,7,11,14,2,-5,10,-5,10,-16,-12,-14,-14,-17,-19,9,-2,20,-6,16,-18,-5,5,-6,-6,19,15,-11,-5,2,18,-11,-8,-16,-4,-20,19,0,15,14,14,-15,0,-7,-6,16,12,18,0,-2,20,8,-7,-6,3,-19,5,13,-3,-20,5,-13,-14,-11,-20,-4,1,5,-17,12,17,12,7,3,-1,1,-10,7,-10,-10,-17,5,17,18,-7,20,-20,17,15,10,0,10,19),
	(9,-5,15,-6,-17,-1,0,9,0,-7,13,18,17,-13,-8,3,6,-1,3,-4,18,17,-6,-15,-4,14,13,-16,11,8,-6,-1,11,15,4,-13,-11,-1,2,0,0,12,-8,-13,4,-7,-15,6,20,7,20,-1,-6,5,-3,8,15,-14,15,11,-16,3,-17,0,-19,16,2,14,1,11,9,-2,-16,2,-18,10,6,-1,-6,-2,1,-13,-4,-12,7,8,-6,19,10,15,10,-19,7,-8,15,-19,7,-13,6,7,-15,-7,-3,8,-15,14,7,-18,-1,20,-15,-6,-10,8,-10,-14,6,-10,-10,-15,19,12,3,3,9,12,2,19),
	(0,4,4,20,5,-10,16,13,2,16,-20,2,3,-19,-19,7,16,3,15,-4,-13,5,-4,18,17,18,-19,13,16,6,0,-8,-2,-6,-10,0,-10,7,12,-13,-13,20,6,0,-9,18,5,2,-18,11,1,7,-2,-16,19,2,-2,-15,14,-2,-6,8,-14,1,-5,10,4,-11,1,19,-3,5,-4,-18,-12,19,9,-14,5,-20,-16,8,12,-13,8,15,14,-17,1,0,0,-7,-14,11,5,12,13,-4,-13,17,-9,-14,18,18,13,8,0,4,18,-1,-14,-17,12,-10,-6,5,14,10,-16,0,13,-7,16,15,3,8,-14,17),
	(4,-8,-12,-5,-12,-3,-14,8,0,18,3,18,-9,15,-20,-12,5,8,19,13,11,-7,-18,-1,9,-5,-19,13,19,-18,12,3,6,-17,8,5,19,16,-6,14,10,12,-12,12,-20,12,16,-11,-17,-3,17,15,-11,-6,16,2,6,20,8,-9,0,8,-2,-12,-18,-20,0,-16,13,0,-17,-12,-13,18,-10,17,-1,-2,-8,-9,8,-18,-8,-9,-17,-14,8,12,1,6,-18,0,-18,-5,0,3,1,-1,-6,-12,-17,7,10,-2,10,16,-19,-2,-8,-11,-16,-9,15,-10,-4,17,-1,16,-1,-2,5,-3,16,15,6,-20,-9,-17),
	(1,19,5,-1,-11,-10,-17,18,8,-1,15,-11,17,14,0,19,0,-15,-7,17,-14,7,-16,18,12,-7,9,7,15,19,-2,1,-4,-3,6,2,8,9,15,-20,12,16,-1,6,19,1,-10,19,13,12,0,0,17,4,-13,-8,7,-1,-14,4,0,8,19,2,10,4,12,1,-9,5,14,11,-13,0,-2,-3,-16,9,0,-13,12,17,7,11,5,-3,-14,14,0,3,20,-18,-16,-14,-9,-5,-2,-2,9,-7,16,13,13,7,16,19,-10,-14,15,3,-21,-3,-14,3,5,10,14,-7,20,-12,-19,13,-12,-14,-10,20,11,-4),
	(-7,-10,-17,-15,14,21,6,-18,13,-12,-7,6,-15,-20,20,11,-21,0,0,-17,-12,-3,5,4,-14,3,12,-11,-1,-6,-10,21,4,20,-18,13,13,-1,-15,-16,6,-4,29,14,0,1,26,-2,6,10,-1,-9,-15,-14,-5,6,-6,-17,-13,-14,-16,14,-16,-5,3,-11,11,-4,-15,13,-6,0,17,-7,25,20,-13,-17,12,4,-17,-12,14,-15,-14,-9,0,-2,4,1,15,7,-5,6,-25,7,-7,19,17,-13,24,-12,16,0,-10,-7,-10,16,-22,-23,-26,11,4,10,12,-11,5,-15,-10,-1,-3,15,14,7,-18,23,2,-5),
	(15,15,-37,-9,-8,30,21,-7,-14,11,16,34,18,-1,38,16,-29,-19,13,-6,-8,-18,-11,4,14,28,-3,3,-8,5,-6,17,-11,-16,20,4,-8,-20,7,5,-9,3,8,6,-20,-19,-2,15,-14,-9,7,-15,8,-24,0,-34,4,-13,-5,2,-3,-6,-6,-20,15,-16,-4,27,-7,6,0,16,-11,-1,16,26,-16,11,-27,-34,-1,-8,-37,-2,6,0,-31,15,4,13,25,-5,33,-1,-4,-3,-10,17,-10,-22,20,2,2,-7,-12,-5,5,21,2,-28,-1,-11,15,-10,-29,30,21,4,0,12,15,-12,30,11,0,31,22,-34),
	(20,25,-10,22,-35,13,10,-17,9,9,-11,0,19,16,0,-1,-35,-19,2,5,-13,-17,-24,0,1,-2,-7,16,-6,23,-11,3,2,16,15,-20,10,0,6,-18,16,15,22,21,-6,-14,36,40,1,23,2,0,2,-31,6,-34,-15,-6,-19,-14,-12,-17,-16,3,5,-17,-11,34,-20,6,2,11,-24,-30,24,2,-31,-6,-2,-29,-19,-31,-11,0,-24,-8,-25,-1,13,-9,28,20,21,9,-38,2,-5,0,5,-12,16,1,-5,5,8,-1,-8,38,-7,-37,-18,-2,28,-3,-10,35,7,-21,-16,1,-12,-1,12,16,36,23,-13,-18),
	(-16,27,-16,-3,-6,22,30,-9,-4,-2,8,3,16,-26,2,-11,-9,16,12,-10,-11,8,4,5,21,-4,6,0,-28,1,-13,33,-6,30,24,-3,0,16,-7,-23,-12,1,13,26,-32,6,21,4,-17,13,-11,6,11,0,-9,-32,16,-15,-2,-4,-12,4,11,-4,11,9,8,24,7,-1,14,-4,-3,-28,27,-3,-12,0,-16,-24,-19,-1,1,0,-5,-31,1,16,3,-14,19,37,8,5,3,16,19,8,25,0,1,0,18,-7,-11,-2,-27,3,-4,-19,0,3,31,9,-35,7,15,-2,-22,-4,1,7,18,35,4,3,1,-22),
	(-9,8,-38,-3,14,15,5,0,-8,23,-1,21,15,-7,12,20,-4,11,1,8,-16,-8,-17,-12,1,3,-9,19,7,-12,-28,2,2,27,20,8,-6,-5,-13,-4,-15,15,21,35,-1,-15,13,18,-24,26,-14,1,-1,-11,-2,-33,-24,-15,-20,-2,3,7,-3,-24,-13,-15,-15,20,-10,-20,19,-12,-14,-25,19,27,2,23,-6,-21,5,-27,-8,3,1,-5,-2,3,15,18,-10,17,19,18,-33,-10,3,37,12,-22,19,20,17,12,17,6,-16,17,-6,-10,-21,-1,25,-7,-34,32,13,2,11,-4,26,0,-4,20,0,18,26,-19),
	(23,52,-4,-3,32,-13,11,-8,9,3,0,44,-9,10,48,12,-17,-19,-11,-10,9,-6,-15,-14,2,4,2,16,-16,20,-41,0,-25,2,-1,7,28,-31,-12,-32,12,27,27,-4,-11,1,23,32,-12,17,6,-14,9,-7,6,-31,-1,2,-16,16,12,7,-10,-17,-23,9,-13,30,-46,-22,32,-15,1,-35,32,-1,-8,-2,2,-6,12,-1,10,-1,0,11,-22,4,26,-8,-3,2,24,-7,-14,22,-1,3,22,0,27,19,-2,-20,-14,-1,-28,19,-27,-8,-21,-11,16,-22,-33,8,24,-22,8,-30,1,-38,19,28,-15,14,9,-17),
	(27,19,-2,-2,33,20,9,-19,5,10,-20,10,5,6,4,21,-18,-6,-3,-12,-27,-5,12,5,24,8,-2,-6,-6,-6,-22,7,-26,7,-1,-18,12,-5,-29,0,-6,2,49,9,-15,-30,26,33,-18,28,25,-18,14,8,-10,-38,-15,-21,0,-4,13,-32,-1,0,15,7,15,15,-46,15,7,1,23,-21,-4,27,-34,9,-26,-3,18,-7,20,1,-16,8,-20,10,21,21,5,5,16,32,-11,-9,8,-10,1,-26,-2,20,6,1,-13,38,-35,14,-6,8,3,-29,4,1,-44,11,33,-21,3,0,8,5,5,7,12,1,3,-15),
	(10,30,-15,2,-10,-10,17,-35,-26,30,6,46,5,-2,1,-2,-16,3,18,-5,-1,-5,18,-13,2,-15,-18,-11,0,26,-38,29,-13,37,-25,7,-13,5,-2,-10,13,8,17,38,-43,-30,10,14,-17,7,-10,-22,23,0,-40,-9,1,-16,-10,3,15,-5,-13,7,-16,0,3,9,-37,-2,26,8,31,-35,27,17,-43,-13,-2,-11,25,-2,5,-22,-7,-16,-13,13,-4,27,4,30,31,36,-26,30,14,18,-7,-21,30,51,12,-4,13,28,-23,17,-5,15,-12,-1,30,-30,-24,32,6,-3,-23,3,3,-13,19,-10,0,32,7,-34),
	(13,31,-40,-13,-1,-8,42,-34,-13,40,-1,48,-8,-27,-1,11,2,13,-8,-20,0,24,5,1,12,8,-31,15,-20,21,-32,0,-2,33,-9,-5,9,-33,-8,-37,18,-8,47,35,-28,-36,37,20,-45,24,9,0,11,-27,-4,-44,-14,11,-18,1,-6,6,-8,-8,3,17,-5,26,-50,-18,4,9,5,-32,9,10,-8,6,-8,-14,10,-6,-7,-17,-18,-7,-8,-12,32,13,-5,-6,-3,29,-40,1,1,13,-1,-8,34,19,13,-19,0,38,-18,5,3,10,-18,14,34,-44,-15,11,21,-22,13,-10,10,-7,21,-16,14,33,49,-24),
	(-26,41,-16,12,-23,-3,-9,-22,11,-3,7,32,10,16,-17,-5,-6,0,-26,-26,6,29,25,2,8,11,1,1,9,14,-5,-16,-4,33,31,4,-21,-10,32,-34,-5,1,10,48,10,24,-4,-2,-8,10,-16,7,-12,13,-6,8,10,10,-2,4,-32,23,30,-2,15,16,15,-15,-19,0,-4,5,-25,-1,15,-3,-1,4,23,8,-20,-11,6,-16,37,4,5,11,7,20,15,-1,-31,30,-27,14,0,-9,-13,22,-25,1,-5,15,40,-12,1,-36,-35,5,20,32,-34,-32,15,-21,-21,-12,-3,-34,13,24,6,40,0,-14,10,-5),
	(-28,55,-39,22,-24,-12,-8,-4,15,16,11,5,2,-14,5,26,7,15,-10,-28,4,-9,-85,7,-17,23,-34,-14,-3,-2,-17,18,-25,41,2,-3,-23,23,-8,-47,22,-9,51,39,-50,7,30,35,-17,-5,14,-28,22,14,-8,-40,12,11,5,20,-2,-6,-8,-4,-1,3,32,5,-1,-7,31,29,8,-2,24,-12,-22,10,-26,-15,-14,-12,-5,-14,40,0,6,-3,-18,21,0,12,29,32,-20,-18,5,-19,29,-2,-16,-13,-21,12,50,0,-23,-16,-19,-19,-17,-17,-15,-45,-15,-1,1,-15,-21,-23,10,9,-1,37,-18,48,-6,-29),
	(-15,16,-29,24,-54,-28,36,-8,10,16,3,6,15,-59,-30,42,2,19,29,8,15,-11,-80,-5,23,-1,-11,12,-37,9,0,-24,39,42,-8,-21,17,-1,-12,-32,-9,-23,52,46,-26,-43,28,17,-22,-35,3,14,3,-18,6,-16,-7,6,-11,-16,21,35,28,-11,-8,-8,-21,19,41,10,9,1,-4,31,-21,6,-25,35,-35,10,5,-15,18,-33,2,-8,-23,0,0,17,-4,18,9,45,-24,0,-9,7,-3,-21,34,11,16,14,0,56,-48,2,-43,3,-47,-19,19,-14,-40,25,42,9,-15,-8,3,23,14,16,32,45,27,-30),
	(-27,15,-18,12,-28,-9,57,-18,-8,40,6,10,-10,-46,-25,22,24,7,20,26,-9,-15,-82,8,6,13,-7,38,-3,-2,0,1,22,37,-13,-12,-6,-10,-3,-6,-24,4,37,20,-28,-26,35,33,-28,-39,22,-6,17,1,-26,-28,-13,19,4,-2,4,9,14,-11,0,-14,0,7,15,-14,-1,10,13,-5,7,-1,5,38,-36,-15,0,0,7,-39,8,0,17,17,-13,-11,-10,1,36,47,-33,0,-9,-2,23,-4,26,-11,23,14,3,35,-41,25,-5,17,-12,3,-1,-31,-17,26,44,2,-18,-6,4,35,25,33,39,41,13,-16),
	(36,43,0,-21,-23,17,14,18,-35,7,-7,27,-15,-6,6,14,-29,6,2,-13,-6,-15,-55,-22,25,-5,1,0,-7,28,-17,27,-45,50,-32,1,-12,-11,-13,-7,-3,33,11,28,-28,24,24,34,-16,21,-16,-9,49,1,-20,-11,37,0,-7,-6,30,-42,-36,-19,-9,7,-12,8,-29,-25,34,-4,57,-18,41,15,-20,-37,9,-56,11,-19,-1,6,-4,8,-19,17,13,22,12,9,30,37,-25,27,9,-5,17,30,16,24,23,-7,10,-2,-40,43,7,-3,-40,-25,34,-11,-38,32,36,-6,13,-18,9,-16,3,6,-2,50,-11,-28),
	(33,40,-24,-12,8,36,6,-17,-29,22,-24,1,0,13,32,12,-39,0,-16,-41,-8,14,-38,-20,-13,18,-14,-18,23,34,-32,38,-19,35,-23,11,2,-46,10,-25,5,51,20,7,-43,-13,44,35,-13,27,-23,-37,34,7,-45,-33,15,-9,-11,4,13,-18,-43,-17,10,1,10,26,-23,0,45,-20,30,-2,51,28,-46,-20,-22,-52,-1,-39,-36,2,5,-18,-20,1,44,-11,39,17,29,4,-13,12,-18,8,37,24,16,11,24,-10,-7,8,-45,52,-20,-7,-25,-23,39,-23,-5,9,35,-18,-16,-19,21,-47,40,17,13,15,-9,-36),
	(40,11,-46,-14,-26,16,23,-11,-40,7,-16,18,-3,22,22,21,-29,9,9,-8,-33,12,-8,-22,18,1,0,-1,11,11,-2,17,-21,50,-18,0,-5,-53,-6,-15,-6,24,15,31,-19,-16,16,30,-23,63,-15,-14,13,-13,-35,-16,24,-17,-19,-19,34,-17,-41,-23,-3,-18,38,18,-18,-15,32,10,52,-15,33,-4,-30,-27,3,-28,-19,-36,-20,4,-14,-9,-15,11,36,0,0,27,38,18,-49,13,5,35,17,-12,15,28,29,-26,0,37,-18,62,-15,-9,-45,6,33,-28,-52,26,25,16,-9,-5,0,-21,35,14,22,27,-3,-11),
	(17,9,-6,-6,-17,38,26,6,-24,14,-22,7,-26,36,40,-5,-13,0,-4,-14,-11,6,-31,-15,-8,31,-22,-7,0,7,-32,17,-41,36,-2,0,0,-11,-6,-24,17,24,35,18,-24,-9,27,20,-44,17,-49,-20,15,6,-19,-16,-2,5,-41,-4,39,-18,-27,-10,-12,6,18,28,-33,-25,27,-10,24,-18,2,4,-44,0,-5,-8,12,-10,-17,-13,-7,2,-10,16,12,8,16,12,38,21,-26,-11,8,26,26,-3,24,40,42,-17,-14,21,-9,14,-19,-20,-9,-1,36,-20,-49,20,32,8,3,9,-8,-46,19,2,-9,31,15,-16),
	(28,38,-12,-7,0,42,12,-12,0,21,-7,30,14,28,21,25,-13,16,0,-20,0,0,-23,-33,-1,33,-7,18,11,20,-11,42,-3,34,-29,-13,20,-5,-3,5,-8,27,30,20,-38,16,31,25,-34,23,-1,-34,25,-9,-3,-28,6,11,-39,11,34,-16,-26,-15,-10,-13,7,24,-8,5,15,-5,46,-31,10,5,-40,-2,-3,-25,-12,-36,-23,-31,-19,-27,-14,9,36,-9,26,-14,25,37,-29,12,8,26,26,-24,0,25,14,-24,-13,14,-3,12,-21,-33,-24,2,12,0,-31,3,28,1,4,0,-7,-43,0,-5,27,26,27,-31),
	(-1,20,0,6,-12,-5,29,5,-7,-1,-17,20,8,24,33,-7,-22,0,-13,-11,2,17,15,-13,-5,19,-36,-4,-2,12,-23,-1,-29,-6,9,-18,0,-19,-6,-16,0,27,29,28,-17,1,0,34,-30,-2,-10,-12,23,-4,7,-2,-17,6,-18,18,2,0,10,-15,12,-10,14,33,-28,-15,19,3,5,-28,-8,1,5,-7,-22,-6,9,-23,-4,-18,8,-30,-20,13,36,-21,29,19,3,10,-34,8,17,14,37,-1,19,20,0,-18,3,-4,-23,33,-16,-34,-33,5,16,13,-35,0,4,-9,-6,13,-11,0,2,4,0,10,0,6),
	(3,0,3,-14,8,-13,-2,18,17,-12,0,11,10,0,0,-2,-4,-17,15,-14,-15,2,20,9,-19,2,9,11,17,8,-4,11,0,-5,-17,-13,-20,10,-13,-19,-16,-4,-18,5,-15,18,-6,-9,10,-20,0,3,16,-16,2,20,3,-5,-4,-11,-6,-3,-19,-2,4,9,3,18,4,-12,18,-1,-8,19,-16,0,-2,5,-12,11,-3,0,19,-16,-19,3,-15,-12,0,3,-14,-4,19,15,3,6,6,1,2,-18,0,-10,-6,-3,1,10,-16,7,13,-9,-19,-14,1,13,5,-3,8,0,1,-16,-5,-10,13,17,10,-19,16,-19),
	(15,-3,-10,12,0,-2,16,20,-9,15,-17,4,-8,-14,1,9,19,-1,6,3,-15,11,-11,6,-20,17,-9,-7,9,-19,-13,-10,-10,-11,5,16,17,-1,-4,11,14,-12,-6,-8,16,19,1,4,19,8,9,16,-12,0,15,-17,7,-6,15,17,-1,-9,-15,-6,12,-8,0,-12,19,4,-10,15,0,-17,-15,-13,0,19,-16,6,4,0,5,-13,-17,-4,4,-13,12,20,11,8,9,13,17,5,-7,-16,5,-2,1,-11,5,-5,13,-14,-12,17,13,-10,0,6,18,3,3,3,-5,7,14,5,4,20,-11,17,-19,-3,3,18),
	(2,-9,8,-6,-17,14,13,-7,-4,3,13,17,15,-7,-16,0,-11,1,-2,-10,7,-14,-19,-1,1,-9,13,-19,-5,-7,-3,20,-15,-11,-6,-18,9,-11,13,-8,-2,-2,-19,17,11,17,-9,-6,-3,0,-20,15,0,3,19,0,12,18,17,4,0,8,7,7,-15,1,-20,14,-12,3,11,17,-19,15,-15,-11,-13,-6,-7,12,-17,-3,-9,2,1,-18,12,15,-9,18,-15,-17,17,16,-19,-1,-16,-15,-7,20,11,4,18,7,9,-20,0,-2,-1,12,18,-14,-20,17,7,-14,13,-9,17,17,-18,-5,-19,13,18,2,13,-11),
	(-12,4,4,18,-19,15,18,-18,0,15,7,-6,19,-8,-4,-12,19,13,13,5,-12,2,6,4,4,2,5,13,4,4,-6,4,-16,0,19,-19,5,-7,11,2,-7,2,-11,-12,-18,16,-6,6,15,-12,9,-2,-12,18,-7,4,9,-3,-18,-17,10,18,-3,11,4,6,-9,-7,-16,-13,13,6,0,14,-2,4,-12,4,-5,-13,2,0,-11,13,0,-11,16,4,-16,-6,-4,20,13,0,19,3,4,16,-11,10,-1,-17,-3,2,0,4,-12,-7,20,7,7,-2,4,-18,-3,-12,-11,2,-2,-16,-14,-8,6,20,-16,-18,14,5),
	(-5,-3,1,-15,-17,16,-16,9,-4,11,-15,-1,-16,1,13,-8,11,-15,-6,10,-1,16,10,-14,3,-9,16,-9,-19,20,-11,9,-15,-18,4,0,2,-18,6,-6,14,-18,0,-18,9,-13,-19,10,-5,5,-14,3,-3,-8,5,-3,-12,13,15,-10,10,2,-4,-20,-15,-7,-11,13,12,0,-19,9,14,20,-14,-8,14,-15,-10,-8,2,0,6,18,0,12,10,-7,-4,1,1,19,0,-9,-12,1,-19,18,-3,19,-15,-7,-11,-12,-20,16,7,-2,-7,1,-11,-14,12,10,5,-11,-12,20,-17,-4,6,8,-15,-15,0,1,18,-18),
	(5,-8,-14,-10,-7,13,-13,-4,18,9,7,-10,11,1,20,-12,-7,9,-6,-12,18,15,0,5,-13,7,0,-9,-14,-4,-15,-9,-18,4,5,10,-7,-3,-2,-5,16,7,-7,-19,-2,-20,0,0,17,13,-19,-9,-16,-5,-16,-18,9,-17,7,-19,-15,-12,16,9,0,-13,-3,2,12,13,-15,4,19,-4,9,-8,3,-15,3,-17,-16,-10,-16,-8,-10,-2,7,8,6,-3,19,11,-13,9,4,6,15,16,-13,-7,18,13,-9,0,0,-11,4,-14,-15,2,-16,-16,2,0,-12,-6,-10,17,10,-14,8,-1,5,-14,10,7,13,12),
	(-15,15,-6,0,-11,-18,19,18,14,5,9,-11,-5,-9,-2,20,-19,-12,-9,0,17,1,2,6,1,13,11,7,1,2,-8,9,3,-9,-11,8,-19,-19,8,9,-18,17,11,-16,-13,0,7,20,-9,0,13,14,17,0,7,-14,16,-7,15,18,12,-8,18,-15,-8,-5,-1,-15,-3,1,18,-11,9,-20,16,-1,-12,13,-12,-17,-5,-17,-3,-8,14,0,1,11,9,0,9,5,-17,20,7,-17,-10,15,17,9,5,0,19,17,16,-10,12,3,-9,-10,16,-5,-5,-3,3,3,-17,4,-5,-2,14,-12,21,13,3,7,4,3),
	(-8,5,-14,26,18,0,4,14,-10,1,14,22,16,1,-7,14,-5,-12,8,-7,8,11,21,28,-1,-27,-31,17,-3,12,-20,-5,0,10,-2,-20,-25,5,-12,-28,12,16,-18,-1,-10,14,-4,-17,-15,-25,24,5,12,-7,8,-28,-16,19,23,18,29,-9,-2,-22,0,10,6,29,8,-9,-16,4,15,-19,-13,15,-35,5,-4,-24,-5,-8,-16,-20,15,-13,7,-12,0,18,-27,28,9,6,15,-11,9,-15,-21,-33,8,-19,27,27,-9,34,-33,-21,-21,3,-16,17,-24,10,-7,36,41,-15,8,4,14,21,-11,5,30,-9,-9,-12),
	(-3,34,5,-12,-18,1,2,18,10,19,11,5,6,-13,-32,0,1,-11,12,15,13,20,-5,-19,20,-12,-32,14,-14,-8,-26,-4,22,1,-23,-3,0,-4,-18,-6,-4,31,26,12,-2,-15,-7,-25,-34,-2,2,11,33,-14,-8,-24,10,-1,25,-16,27,-18,-11,-22,5,18,-4,2,-6,5,22,18,24,-18,6,-12,-20,13,-18,-11,9,6,2,7,4,1,7,-9,-7,10,14,7,11,3,-3,-12,-7,-9,2,-32,-13,-25,-9,13,-9,35,-30,11,2,2,11,3,-12,-22,-28,18,13,18,-19,-3,14,7,-10,19,4,-3,-15,-8),
	(5,3,8,11,-4,14,17,10,1,-16,0,-5,-4,14,26,12,10,-15,8,4,-20,-8,7,12,-15,24,8,-8,15,-11,20,8,-9,13,-14,-13,13,6,5,-17,10,-11,40,40,-13,-19,24,25,-30,0,7,12,-1,4,-30,-1,-1,14,4,5,-2,15,-10,-3,-3,-13,-6,9,5,0,8,-4,-1,-1,26,17,-9,-20,-18,10,21,18,-17,-2,8,18,17,15,16,-4,-7,-12,-10,2,-9,-5,-19,26,18,-1,10,-1,13,17,-6,5,-9,-10,-22,21,-20,-16,1,-19,-5,18,7,-13,8,-29,-13,1,-6,-6,11,-17,27,-23),
	(13,30,-34,-14,0,5,14,-20,5,8,-1,32,20,4,28,5,-8,0,15,0,0,-36,-33,16,-19,22,-2,-16,11,10,8,22,-15,-6,14,-29,17,-2,-31,-11,0,11,29,8,-7,1,45,11,-26,28,-15,-24,-16,-36,-14,-15,6,-15,-32,-16,-7,-22,-11,-26,-19,-14,10,28,-34,-15,29,-14,26,-26,23,6,4,10,-13,-9,7,-24,-4,0,0,-6,-35,26,-1,7,24,-14,31,3,-37,0,12,28,13,-1,31,16,24,-5,-11,26,-30,18,-30,-19,-38,-13,32,-10,-13,7,2,8,-9,-15,0,-3,12,55,15,18,15,0),
	(10,13,-36,14,-8,-10,29,-21,-30,36,0,35,-6,4,18,14,-21,-5,10,-5,7,21,-28,23,-6,16,-12,-15,17,-6,-4,26,-12,-6,-6,-18,-15,-5,-9,-20,-12,6,7,16,-42,0,35,1,-20,-4,-20,-37,22,-33,-21,-28,5,-20,-2,-12,9,9,-20,-24,-18,-22,10,14,-34,-23,13,-20,12,-34,39,14,-32,8,-34,-9,-2,-33,4,-2,-17,1,-24,6,24,-2,9,12,35,20,-17,-5,-21,20,1,-20,19,25,-1,0,17,29,-25,25,-15,-16,-36,-17,6,-15,-18,23,20,-28,-9,3,-7,18,33,29,31,8,19,-32),
	(-6,12,-9,0,17,38,16,-13,3,0,20,2,0,11,18,34,-14,-17,1,-24,-7,1,-48,-19,3,46,-6,27,41,22,-11,41,-11,8,49,-32,26,3,-23,-22,-5,-10,45,39,-8,-23,24,33,-33,13,-18,-22,15,-38,5,-45,-13,-4,-20,-16,3,13,6,-24,-6,-9,22,37,1,-32,12,8,15,-40,1,18,-12,0,0,2,8,1,5,-22,-37,4,-20,21,-7,-24,5,-17,48,25,-22,-2,15,39,-15,-2,12,19,24,1,1,21,-33,14,0,-2,-28,-12,20,-38,-49,19,25,-27,-13,0,8,0,12,20,23,0,30,-33),
	(-4,0,-49,16,41,37,15,5,4,-5,20,-5,-16,2,44,42,5,-11,-2,13,-20,-15,-12,3,-21,66,-46,14,24,-13,31,19,1,-10,60,-11,8,3,-18,-37,3,-22,42,54,-2,-22,10,32,-58,30,2,-4,-17,-11,-5,-30,-13,-35,-42,-6,-27,30,-11,-25,2,-27,-11,0,4,-5,52,26,10,11,2,40,9,9,18,-13,-26,5,60,-6,-17,-27,-17,12,-1,5,-20,-20,7,7,-28,17,-2,19,-48,6,23,-4,0,-7,-33,47,-27,4,-16,-30,-23,-18,18,-17,-26,22,7,16,-26,35,45,11,27,39,49,-14,35,-7),
	(0,19,-34,1,14,18,49,2,20,33,16,-6,10,-13,23,42,14,-1,28,-14,-31,-37,-16,-22,-8,60,-41,0,33,-10,0,19,19,-16,33,-14,24,7,-54,-18,-2,-24,39,45,-8,-54,39,25,-69,3,-12,0,-1,-2,5,-7,-41,-25,-39,-14,-7,15,0,-17,-37,-55,-12,6,1,-5,37,6,-2,20,1,36,1,5,-24,-10,-42,0,35,-37,-14,-9,-23,-7,-8,11,0,-18,28,31,-38,-4,32,34,-29,-34,59,21,16,14,-29,26,-48,40,-11,-16,-20,-30,5,-19,-44,31,20,-10,-46,43,28,9,57,30,18,6,57,-24),
	(1,45,-38,11,4,26,57,-13,20,48,11,31,16,7,32,24,21,-8,11,20,-52,-18,-56,-29,-34,50,-14,39,8,7,8,1,19,13,-8,-10,24,-8,-27,-25,-48,-8,85,81,1,-34,44,12,-61,-5,23,0,-19,-24,0,-6,-41,-9,-30,-4,5,22,-19,-26,-12,-53,-13,28,0,-15,77,20,-31,7,19,43,-23,11,6,3,-29,-4,13,-35,-10,-30,-16,22,25,5,5,13,26,14,-67,-25,0,52,-28,-19,10,4,-11,1,4,62,-21,47,-38,-12,-31,-14,12,-8,-82,44,53,-29,-8,12,5,-16,58,-8,42,-2,29,-32),
	(-5,29,-20,6,-44,19,40,6,-12,9,0,0,20,-20,44,51,28,17,23,5,-30,-17,-46,-12,-39,33,-42,20,11,6,17,30,1,-9,24,-2,4,4,-7,-17,-13,-26,34,37,-40,-37,32,31,-26,-1,-8,-10,-6,-19,13,-39,-15,17,-28,-12,-2,31,20,-34,-15,-44,-23,29,-14,-34,42,42,0,5,3,32,4,28,-1,-13,-24,15,16,-40,10,7,-33,40,11,-4,-1,21,23,31,-47,-40,-3,12,-44,-27,28,15,21,-6,2,47,-50,19,-61,-12,-67,-35,30,3,-85,26,12,-13,-52,9,-2,-3,39,25,18,31,29,-39),
	(-16,32,-31,31,-45,19,-2,-5,-10,-19,10,-22,-15,-34,36,-5,61,-8,-17,8,19,-12,-1,-26,-44,11,-36,12,42,-6,-11,44,-28,32,20,-51,-16,-4,1,-30,11,-19,48,38,-40,0,0,76,-56,-1,-17,-17,-17,2,21,-13,-12,-6,-49,14,-25,21,34,0,-8,-39,-35,1,-27,-26,55,20,-53,-2,24,1,-31,24,-18,-11,-32,-38,12,-47,25,5,-6,10,-5,-1,42,-25,-2,45,-49,17,-19,-13,-28,15,-8,43,-17,21,-5,4,-58,9,-44,4,-21,-32,-16,-40,-71,18,-13,-4,-69,10,2,11,33,43,2,4,-5,-12),
	(12,14,-46,10,-61,39,21,-6,-3,-27,23,-24,-23,-52,47,17,34,-10,-6,14,-11,-5,11,-15,-35,45,-31,0,19,-24,28,32,-20,-7,34,-46,-11,-12,-18,0,26,1,60,82,-22,-18,33,35,-23,0,-3,-11,-61,-11,7,2,8,-13,-35,-5,-42,32,29,8,-8,-54,-65,-1,-53,-15,34,8,-46,-21,41,8,30,7,25,-16,0,-28,27,-59,11,7,-26,37,-8,-4,18,-23,12,16,-57,57,0,-17,-19,-17,-1,44,-17,4,-12,19,-55,49,-45,-20,-22,-12,22,-22,-32,22,3,-5,-60,-18,-11,17,57,10,40,21,33,-21),
	(-7,18,-43,22,-92,9,3,-20,3,11,10,-6,6,-38,62,34,33,-4,-21,-28,2,-25,-20,-7,-42,19,-4,-7,48,-31,37,44,-41,24,27,3,-32,11,-43,-4,41,27,11,71,-57,32,11,45,-38,-17,7,-34,-22,2,5,0,17,-7,-72,-16,-24,28,22,-15,5,-45,-50,19,-13,-8,67,17,-62,-52,50,0,1,16,24,-17,0,-4,13,-55,6,-27,-32,38,-4,41,20,-36,-18,31,-87,52,-35,22,19,-26,-13,28,5,25,10,13,-52,11,-41,-8,-28,-21,11,-23,-45,-7,5,-17,-63,-5,1,8,48,-38,17,20,-7,-43),
	(-20,14,-33,9,-62,-4,-1,-36,-14,25,-14,14,33,-64,20,29,18,29,-25,-21,-5,-20,-34,-12,-5,21,-12,-11,36,23,5,44,-43,38,42,0,11,30,-37,-4,55,43,10,6,-42,25,26,24,-38,-19,-12,-31,10,14,17,-9,-8,-27,-61,-9,20,20,8,-39,-19,-51,-42,18,-22,-2,46,24,-32,-44,29,-20,-10,-7,-23,-32,-21,-37,10,-68,13,-31,-12,37,2,-6,0,-29,-9,41,-57,39,-22,-7,30,-13,-10,-9,-10,19,-4,-7,-12,2,-20,-16,-38,0,10,-16,-14,18,6,2,-16,-4,5,12,2,-46,15,46,1,-33),
	(21,9,8,32,-42,7,-9,-35,-36,-3,-6,30,11,-53,16,4,-15,-3,-15,10,17,-19,-38,-6,-12,48,-2,-28,6,37,9,43,-4,25,41,-18,25,10,-22,-4,15,21,10,9,-12,11,-1,36,-9,-22,-27,-36,5,0,-4,-7,-10,-28,-44,17,9,24,-7,-33,-6,-47,0,29,21,-26,35,7,0,-26,33,4,21,-11,-22,-19,-6,-17,-26,-41,7,-38,31,33,26,4,21,-27,-6,-12,-45,29,-25,20,50,-9,-4,-14,12,19,-11,-6,-1,11,-2,-25,-9,-23,-6,-13,0,4,-5,19,-24,-2,0,-19,39,-7,-7,44,18,-42),
	(9,0,-19,0,5,-4,16,-12,-34,0,-16,-9,-11,-51,-3,27,-13,-2,3,-2,20,-9,-27,2,16,38,-4,-6,-32,48,13,22,3,17,44,-5,32,18,-10,13,16,45,-2,-13,0,-8,-1,68,-22,-16,-44,-26,-2,14,14,-8,17,-29,-21,14,34,7,5,-16,-27,-16,12,12,24,0,-2,15,23,-54,47,13,23,-27,16,-18,-38,9,-44,-47,13,-18,20,11,2,6,-12,17,18,-12,-25,49,-26,8,4,-22,28,7,7,15,-8,2,-1,5,-17,-12,0,19,18,6,-10,-19,16,8,17,-4,21,2,3,64,-15,22,40,-41),
	(5,-1,-7,-19,9,3,-24,-3,-38,-15,-59,7,-10,-37,11,-17,-8,-9,-42,-28,-24,13,8,-32,-4,-8,-8,-49,-12,8,2,4,-41,55,11,21,-3,0,3,0,1,41,-24,9,-12,10,-6,57,-11,17,-9,-7,28,13,2,-19,17,-20,-28,0,26,-7,0,-1,3,13,10,30,-28,-19,2,7,45,-27,29,32,-19,-9,-9,-32,5,-33,-1,-24,2,-24,39,42,9,-16,19,-10,10,2,-82,40,-3,0,56,-40,3,-19,14,12,-6,-36,-11,0,-2,10,-32,0,15,8,-22,-4,-2,17,20,33,-7,24,8,34,14,27,-2,-36),
	(49,4,-17,16,13,-7,21,4,-43,19,-49,11,-21,-37,-21,3,12,-9,-56,-21,-19,15,-2,-29,-23,30,-17,-15,20,14,14,0,-4,43,10,2,18,8,-19,2,29,37,-6,35,-23,24,11,70,-26,29,-6,-30,29,20,-19,-50,12,-17,-39,-19,20,-19,-19,-9,-15,-6,-23,22,-44,0,27,-6,21,-23,11,25,7,-22,9,-19,6,-16,9,-14,10,10,12,21,14,-17,25,17,13,-6,-39,60,-20,0,28,-16,22,10,37,-16,-26,20,-29,42,-16,-24,-46,0,-1,-1,-24,25,26,8,5,25,3,-14,-9,27,23,32,-7,-39),
	(52,-3,-20,-10,17,0,59,5,-30,34,-40,16,-11,-22,9,13,6,-9,-9,-8,-35,1,0,-49,-18,13,4,-23,12,7,6,27,-13,13,1,-28,-7,-3,-33,-35,8,30,-23,40,-45,16,42,78,-38,44,0,-24,18,-5,-18,-36,12,-34,-47,-9,-1,-32,-10,6,-41,-15,-29,34,-42,-4,4,17,51,-7,26,27,-17,-17,7,2,8,-3,7,-9,10,0,9,2,38,3,-1,25,22,4,-27,0,-3,47,42,-15,39,30,43,8,-13,40,-33,33,-25,1,-35,23,36,-46,-40,43,16,0,-11,7,6,-20,0,56,30,26,33,-22),
	(33,21,-19,4,33,28,16,17,-13,20,1,19,-15,-15,0,-13,-17,-15,-16,-16,-17,14,3,-33,-2,22,-10,-23,25,-5,-23,38,-38,52,-16,-12,2,-30,-5,-16,12,26,19,35,-24,3,44,50,-1,64,-12,-42,13,25,-2,-18,3,-13,-12,-8,24,-28,-39,-7,-20,20,-30,17,-14,-2,8,4,34,8,31,9,-36,-15,20,-32,6,-44,5,-28,-20,24,10,16,52,7,35,31,43,34,-40,18,-10,46,23,-11,6,39,35,-25,-10,6,-32,30,-11,-7,-20,6,20,-32,-27,19,37,-3,4,-10,11,0,27,46,12,10,32,-34),
	(32,17,-13,-4,-10,12,14,15,-18,24,20,23,-22,-15,0,25,-20,-17,14,-1,-19,-36,-37,-30,-12,8,-33,5,17,-5,-1,9,-28,38,5,-21,-15,4,7,-13,2,25,0,30,-22,18,2,54,-45,20,-32,-10,42,28,-20,-52,1,-22,-24,-12,20,-23,-20,1,-1,-1,2,24,-16,-16,-9,0,30,-18,22,-5,-22,-9,12,-33,-23,-25,-20,-25,-26,-25,5,5,9,0,24,14,45,20,-44,5,0,28,44,-21,19,4,34,-27,3,35,-18,19,-27,0,-32,3,28,1,-57,24,5,12,-16,24,14,-12,15,22,25,5,22,-33),
	(19,0,-25,-9,-21,0,31,-1,9,-6,-5,-9,7,-20,17,28,19,8,28,12,-12,-17,-5,-31,-19,9,-27,15,4,18,3,-3,-7,3,24,-24,13,15,-5,-11,-15,11,14,2,-26,-10,4,-19,-34,2,-11,-3,-7,30,-5,-38,-35,-21,-42,-8,-14,-3,8,3,20,-21,-4,-1,0,7,-2,24,-9,3,-12,-1,0,13,-8,8,-8,-23,16,-21,9,-5,-7,-1,-3,-1,-17,14,-17,14,-24,13,24,4,-15,-19,34,-12,12,3,-6,19,-22,1,10,9,-34,14,17,-18,24,39,17,-9,1,7,0,-10,13,33,-6,1,35,-11),
	(-20,-17,-23,23,10,-7,31,25,30,-9,32,-12,25,-7,14,31,33,12,4,19,1,-5,-8,7,-22,24,-8,12,22,-2,-1,14,24,7,2,11,8,1,3,-20,-4,-18,27,28,0,21,-21,9,4,22,25,-3,-9,14,-11,-24,-23,17,-11,-15,-5,13,0,-17,-10,-28,-4,-15,23,8,18,10,6,-18,-1,-2,17,-14,-4,-10,4,20,-5,-21,18,-6,7,-21,2,-23,10,-20,-12,-5,0,2,11,-8,-16,8,11,-9,17,4,6,17,5,19,-17,15,-36,7,8,-17,21,18,-8,17,4,9,-12,1,12,-14,-8,0,21,-10),
	(-3,13,1,18,-6,0,2,-11,6,14,-12,12,6,4,12,7,4,-9,10,-13,-8,-18,0,-20,8,5,0,-11,13,-15,-8,-18,4,3,4,2,6,20,-13,16,-14,-10,-5,-12,-16,4,18,19,-5,2,7,-7,-17,4,-2,-13,0,-11,0,-6,-16,-15,4,0,18,-5,-17,8,12,19,-3,-16,8,16,-7,1,-4,-19,14,-7,-4,-14,-18,8,-1,-14,15,10,5,-2,3,-4,-5,-16,-11,-18,-11,8,11,-1,-8,-1,1,-18,-9,-19,5,18,11,14,-12,-10,-2,5,-9,5,0,6,-7,-8,2,-12,3,17,-7,9,-18,-20),
	(10,-16,8,19,9,14,-12,3,5,9,-15,-20,18,14,-6,-18,9,-14,-9,18,17,3,9,4,-11,17,4,-6,-2,13,-18,0,2,17,-2,3,18,-20,-19,-11,-9,-7,-13,15,4,10,-10,-1,-4,19,-11,-5,17,-7,3,-3,7,-20,8,5,-16,-3,-2,4,20,-13,-3,-15,6,2,-18,6,-12,-11,1,20,9,2,-3,-7,9,4,5,-2,-3,20,2,-20,4,6,10,-1,0,-14,-6,-7,15,11,-6,-19,-4,-5,-7,15,0,3,-11,-5,19,19,-20,11,6,-19,-5,-3,-16,-4,-18,-1,-10,-4,6,-19,20,15,-5,17),
	(16,16,-7,-12,-13,5,-14,15,2,13,1,14,18,13,0,3,-12,2,-2,0,-4,-17,11,17,-15,-9,-18,8,-12,19,0,0,15,-7,-7,-5,-3,-1,-6,-8,11,20,15,4,14,-9,-3,1,6,-1,-15,17,2,-5,0,-6,-5,12,-1,-5,-2,6,-19,15,-19,-7,17,13,-14,19,-18,4,7,-9,7,11,-13,-10,11,-15,7,17,-15,0,-3,-17,-7,-15,0,0,-10,-2,7,16,-8,15,-16,-12,-5,-7,9,-3,-12,-5,-4,-17,11,8,-4,20,14,-12,-3,20,-7,19,-4,8,-5,-7,-18,18,-7,-11,18,-20,3,17),
	(13,-18,-14,-14,16,5,15,6,11,-6,-5,-18,-5,-4,-14,-1,-7,10,-17,-8,-11,0,11,8,10,-8,5,8,-11,-11,0,-9,4,-10,4,-2,8,1,-12,12,-9,6,19,-6,-13,18,20,-8,17,-9,0,5,-16,18,-8,10,-15,2,-19,-7,0,7,7,1,-4,15,-18,-18,-14,5,7,-15,14,-3,0,9,16,9,0,-9,-14,6,19,7,-19,-5,7,7,-2,-12,0,3,-7,-12,16,8,-18,-14,-19,12,11,1,6,1,-9,-19,1,-2,-5,-9,-8,-14,-17,19,-8,-2,2,-5,12,-10,-14,-19,19,7,-9,13,17,17),
	(-24,19,-22,27,29,-16,-22,6,18,1,37,-1,23,15,18,-15,-30,27,17,-6,13,0,1,28,5,17,18,17,13,19,40,-33,-7,11,40,6,-7,36,-1,11,18,17,-4,29,-36,46,-41,1,-43,-7,0,-40,-1,5,31,6,-17,-15,-13,7,-38,40,5,5,12,-27,-13,-26,8,4,32,28,-43,28,15,-32,-21,7,6,-34,15,-18,18,19,25,-4,-16,-14,-18,37,33,-19,-16,30,0,-25,13,0,-14,-17,-27,5,-18,20,30,-13,5,-6,13,5,34,10,-4,-33,13,-10,-31,20,29,39,4,-7,9,1,-38,-21,-9,39),
	(13,-3,-19,3,-19,-13,24,3,4,6,-8,-18,7,13,-23,-10,-33,18,25,10,22,-3,-6,-3,-7,-1,2,0,-4,-8,-24,28,-3,39,10,28,5,-15,-38,-30,-4,36,37,0,-17,-15,37,15,-9,-27,18,-30,35,-9,9,-10,-33,-5,17,0,23,7,-1,-23,20,-9,28,26,15,11,14,9,40,-15,11,6,-39,16,-20,-43,-29,-28,-14,9,-13,2,3,6,20,15,-10,27,50,22,0,13,-23,14,-3,-24,22,-22,26,28,-6,10,-24,2,-20,-10,-25,-13,-15,-1,-48,32,7,11,-24,15,6,-9,30,-5,5,21,-15,-17),
	(37,-6,-3,-26,-16,-25,-5,-13,-11,-7,6,-7,21,9,-23,-35,-26,11,7,-14,-3,10,-45,9,32,-2,-18,-23,-21,3,6,0,-3,24,22,-16,34,-4,-3,24,-14,8,-5,5,2,0,12,16,12,-28,-41,-17,24,-14,-5,-19,-10,-13,-19,-4,35,2,-13,-37,-4,35,45,-6,-30,12,-29,-23,39,6,41,6,34,22,-7,-22,14,10,-35,-4,8,-18,0,50,-1,27,16,-20,38,-3,-31,18,3,15,42,-43,34,-13,0,5,4,-14,3,26,16,-6,1,-22,-9,-7,-25,-32,6,-4,-12,12,51,2,19,-18,-25,20,9,8),
	(-24,23,-13,-23,19,-9,-13,24,14,5,-16,-6,-2,-26,27,-19,23,-39,6,12,-27,-3,-31,-13,0,30,-39,-12,20,20,-33,1,20,-18,1,-11,11,-22,6,13,-3,-15,0,9,28,-5,41,-1,-2,17,13,-29,-3,-2,9,-37,8,18,-36,2,31,9,-21,-15,-32,-26,1,32,-30,-14,11,23,1,-19,30,11,6,14,23,-7,13,20,-5,-15,-2,-8,-37,29,32,18,-28,3,12,-3,-36,11,13,14,15,-16,18,0,32,-17,-17,11,-24,18,-26,2,-40,0,17,3,-13,-3,13,-16,-22,17,-4,-16,-3,8,6,-13,-10,-34),
	(-31,4,-13,16,-11,23,-1,-3,0,3,3,3,0,-8,48,8,6,-6,10,-8,-28,-21,-45,-19,-16,25,-29,-11,43,7,3,35,-2,-17,-20,-1,-26,-25,4,14,5,-32,35,2,-20,-24,48,0,6,31,-28,-5,-31,-28,10,-29,-17,6,-48,-12,-9,4,9,0,-13,-38,7,38,-18,-3,44,7,-16,-11,40,14,-29,22,1,-29,-15,0,0,-31,0,-39,-29,13,32,-13,-20,14,27,18,-19,-19,13,31,-1,-17,-1,23,13,-18,-14,12,-31,17,-21,-13,-40,-2,42,-12,-35,19,49,-2,2,-5,-4,5,8,1,6,-2,-18,-26),
	(-1,29,-52,-5,-18,-2,-20,-1,4,37,-11,0,7,22,32,-4,5,-40,-9,13,-17,-34,-20,-10,1,7,-36,21,11,20,-16,37,11,0,-30,-11,-17,8,-2,3,-19,-26,23,11,1,-16,42,-3,-13,28,-11,-8,-10,18,7,-34,-9,-22,-15,-16,28,10,-12,6,-1,-14,14,15,4,-33,48,-7,7,-13,40,9,-26,39,-2,-19,-6,-11,24,-13,5,-42,-39,45,43,2,12,0,6,19,-62,-16,26,42,-22,0,10,-16,28,12,-10,-12,-46,4,-43,0,-28,-18,14,3,-5,12,37,0,-8,36,21,-21,-9,0,18,-9,8,-57),
	(-7,48,-57,16,-10,9,2,56,-31,6,10,-3,8,-4,2,14,0,-26,-9,24,-38,-20,-26,-25,-22,18,-39,39,0,-18,7,23,46,-20,-14,-25,-1,-6,-34,-15,-7,-38,18,-2,17,-48,51,-12,8,9,6,-13,-11,15,22,-35,-15,2,-9,0,11,14,27,-26,-36,-32,-50,35,22,-21,37,15,4,-6,31,36,-18,31,-31,-9,-22,8,15,-46,28,-47,-28,12,13,26,-23,26,18,-11,-77,-12,36,50,-47,3,4,15,19,6,-43,-6,-48,28,-27,-6,-80,-22,31,31,-56,43,66,14,-8,36,-10,-30,-30,-28,-23,13,-22,-32),
	(5,29,-56,36,-21,-3,24,15,-1,-7,20,-9,3,7,8,4,9,26,23,30,-41,-3,-24,0,-27,43,-49,25,0,-17,13,12,51,-16,10,-53,34,17,-35,-28,18,-26,12,23,-7,-31,23,10,-38,29,-22,-25,0,59,16,-34,-8,-20,-15,15,21,28,30,-35,-21,-35,-28,18,-1,-14,55,23,-5,-21,-4,39,-2,34,-45,-25,-15,8,-7,-25,-16,-51,-40,3,-15,0,-24,2,34,3,-66,7,6,47,-39,-23,13,0,17,4,-10,18,-70,38,-38,-3,-45,-32,27,-18,-63,43,38,24,-41,61,41,14,15,-9,30,-9,24,-34),
	(-27,3,-51,25,0,19,4,33,7,6,11,26,-1,-16,-3,27,14,16,-6,13,-71,3,-33,-28,-14,28,-60,19,13,-40,-20,-6,45,-18,-4,-33,-3,25,-47,-9,13,-26,-1,-18,-7,-12,29,0,10,23,-1,-21,0,31,17,-42,-11,24,-26,-20,0,20,24,-43,-37,-35,-27,8,-35,-1,12,28,6,-5,9,47,-4,31,-23,4,-53,31,17,-13,11,-28,-7,4,-17,9,-38,-5,11,-7,-51,-4,24,39,-39,-6,1,11,-9,0,-24,7,-41,18,-48,-31,-59,-30,-2,-3,-89,15,48,13,-33,29,29,-21,8,-2,-4,-24,-6,-47),
	(-4,15,-49,25,-18,13,27,21,20,13,-14,-7,-12,-30,4,12,1,10,-11,41,-75,-12,3,-25,-31,20,-48,10,29,-11,-18,-8,56,-37,8,-23,7,8,-3,-11,-6,-50,-9,-12,44,-27,43,-13,-14,18,-1,16,-31,8,35,-27,-20,7,-17,18,31,24,2,-14,-46,-44,-21,16,-36,-31,20,10,-8,19,-12,31,1,44,-12,-5,-24,38,18,-2,12,-29,-42,28,15,18,-29,13,52,-25,-59,0,15,31,-2,-29,25,37,-4,0,-53,16,-76,10,-37,7,-52,-11,12,-16,-73,27,29,20,-30,30,18,-1,13,-55,13,-35,31,-35),
	(-21,59,-54,30,-65,23,3,35,-12,17,-1,9,-17,-11,26,14,2,23,-8,6,-25,-25,-6,-15,-8,13,-44,13,19,-7,-12,34,15,-25,20,-46,18,9,20,12,26,-31,3,3,19,-6,35,1,-18,-1,11,7,-7,8,9,-38,-8,9,-24,-5,7,48,30,-37,-18,-15,-14,38,-11,-28,36,45,6,5,15,26,9,34,-25,-31,-46,-8,15,-26,21,-20,-28,15,-19,-9,25,-8,24,-8,-65,2,22,21,-13,-2,0,44,-10,21,-22,18,-88,35,-42,-19,-43,-14,30,21,-88,14,42,22,-32,51,-11,0,0,-42,-13,-2,13,-46),
	(9,27,-73,20,-90,-10,27,21,-4,48,-24,6,-14,-65,2,34,-27,32,16,15,-47,-19,20,-22,-28,-3,-13,-5,-16,-31,-2,5,2,23,-12,-28,-10,14,-12,-13,37,-49,-15,-4,-12,-15,26,31,-3,3,27,-26,18,-35,3,-52,-4,15,2,-1,-1,17,27,-31,-45,-18,-25,31,-45,-13,31,20,-31,21,20,-8,-18,19,-10,-33,-44,2,-30,-82,5,-56,-51,12,-12,-7,28,11,18,46,-61,31,-12,-11,-6,15,28,27,-14,12,-10,38,-78,40,-62,-27,-26,-1,-8,9,-98,53,16,0,-65,44,-6,-14,-12,-17,-32,28,-14,-33),
	(-12,23,-41,20,-121,-15,20,-17,-13,50,-25,-24,-66,-87,28,12,35,15,-26,36,-55,-9,13,-20,-28,7,-30,-15,-36,-57,4,27,27,0,-4,-17,-29,-17,2,26,33,-22,-17,8,-7,4,-4,2,1,7,23,16,34,-50,13,-64,-9,19,0,6,27,52,57,-38,-77,-24,-26,24,-50,-6,-12,1,-70,0,19,2,-10,49,-11,10,-16,7,9,-72,19,-1,-37,-15,26,-7,35,0,23,19,-52,48,-11,-11,-1,15,-2,-3,13,11,-66,15,-78,45,-58,-19,-28,-6,28,12,-76,36,23,0,-37,7,-7,-15,6,-22,2,9,-20,-38),
	(-31,30,-57,3,-110,12,27,-31,2,14,-44,-30,-50,-84,-28,2,13,11,-18,13,-50,-3,44,-27,-21,2,-17,-18,-10,-36,23,20,5,9,0,-15,-30,11,-9,8,29,-9,-27,-11,11,18,-25,28,2,-19,-3,-21,4,-28,0,-33,-1,10,13,6,43,41,13,-56,-60,0,-21,20,-33,19,9,0,-65,-29,36,-2,-25,34,-37,5,-13,-5,2,-56,2,-24,11,0,12,7,-8,0,27,15,-47,32,3,23,11,9,-4,-2,-9,10,-37,-5,-29,52,-32,-26,-20,8,25,29,-15,9,-1,27,-21,12,-19,16,-7,-33,-16,30,-9,-14),
	(9,22,-30,14,-65,-3,2,-35,16,49,-29,-16,-21,-69,-15,0,27,29,-20,26,-29,-1,35,-41,-35,24,-11,-1,8,9,18,28,7,-2,-4,-16,3,-1,-37,-3,29,8,-36,7,-15,14,-10,15,-2,-30,14,4,-8,-29,13,-35,-6,-9,-3,1,28,30,45,-80,-57,-35,3,17,-16,-18,7,22,-44,-51,19,-21,-6,16,-49,11,-44,-27,13,-69,37,-19,-31,7,14,12,11,-4,-41,1,-39,34,-10,18,3,-26,12,-19,39,19,-47,2,-31,11,-30,-5,-22,3,5,13,-12,47,19,-19,-60,-26,-33,2,-2,-38,-16,14,10,-4),
	(-13,17,15,8,-2,-10,15,-57,-2,32,-47,-20,-12,-65,17,-7,-19,-1,-26,14,-14,17,-5,-47,-1,-12,-36,-25,-16,36,17,5,-12,46,1,-2,30,7,-43,10,-8,13,-20,-27,-3,21,-23,2,3,-24,32,10,6,-41,2,-44,-25,5,-5,-16,15,62,12,-53,-75,-4,26,23,-2,11,21,30,23,-64,-1,-7,-9,8,-47,-9,-49,2,-17,-73,18,-35,2,24,0,-23,-3,4,-27,19,-13,28,4,14,7,11,-2,-10,19,0,-23,0,-7,-9,-14,-32,-12,-15,-18,0,-12,29,-6,-22,-14,-14,-30,-31,-3,-7,-15,34,11,-4),
	(-5,13,31,12,5,11,-18,-28,-5,-15,-31,-12,-21,-55,-6,7,-10,15,23,22,-3,-13,-35,-33,-7,12,14,-49,-12,5,20,32,9,42,-20,25,18,2,-43,-4,11,21,-36,-25,12,0,-13,19,0,-17,-26,-20,18,-9,-20,-30,-23,-20,-26,-13,41,43,-13,-44,-66,23,41,18,19,1,19,19,6,-55,19,5,-10,3,-50,-21,-53,9,-41,-27,1,-70,-10,29,19,-36,29,34,5,6,-23,48,-40,7,38,-28,7,14,32,18,-36,-10,15,-2,2,-38,6,28,24,26,-3,11,20,-39,-31,-20,20,-29,-45,2,-52,44,3,7),
	(-3,4,7,-23,22,9,-7,7,-38,5,2,14,13,-38,-13,7,-9,5,24,-13,-18,20,-29,-25,5,-1,9,-18,-31,13,-6,27,7,40,-16,-10,17,-4,-21,-6,-9,3,-9,-12,8,7,-6,40,26,-5,-33,-14,6,-17,-4,-29,-18,3,-24,4,4,27,-19,-45,-25,-8,4,30,8,6,17,28,15,-58,29,16,17,-16,-28,-33,-9,1,-31,-9,-4,-40,4,50,1,19,3,17,-31,-31,-9,11,-30,17,26,-15,-6,-13,19,26,-46,-33,-3,-16,-8,-19,-26,18,0,9,23,-3,22,-17,-16,11,33,-38,-35,2,-12,31,0,8),
	(-5,-5,-3,-12,10,-23,-36,-18,-14,0,-34,1,-9,-10,-26,-26,-11,-2,21,0,-33,38,-39,-54,-1,-28,11,-21,5,2,-8,25,13,2,-2,32,1,26,-7,28,16,-15,3,-23,28,5,-7,-11,53,2,5,-8,-23,-4,2,-31,-12,-10,-26,12,55,15,-11,-43,-54,22,15,-11,-34,23,-10,16,26,-46,34,15,-18,4,-9,-22,-17,11,-46,-17,-2,-23,12,23,-7,7,-8,1,-34,-25,-12,-8,-5,21,20,27,0,3,41,4,-63,-33,-24,-10,-21,0,-33,0,-14,47,0,-4,17,-13,-39,19,32,-21,-19,-34,-33,36,-15,23),
	(12,-21,4,3,7,-4,4,-26,-14,-25,-34,-12,-12,-21,6,-16,-22,-11,7,-11,-28,35,-12,-43,-3,9,26,-48,-8,5,-5,-17,10,53,0,3,19,-12,-14,10,22,35,4,-26,27,3,3,61,12,-1,-41,-15,-11,-3,-8,-44,43,-19,-22,0,17,-10,-11,-39,-68,15,13,19,-1,48,-12,-12,35,-53,48,8,40,-18,-2,-6,22,15,-5,-34,-9,-24,22,2,11,1,-19,8,7,-27,0,17,-17,27,29,31,18,41,1,-11,-8,-12,-26,-33,-25,18,9,-18,1,4,22,-15,9,9,-18,-21,8,12,-18,-40,2,42,5,4),
	(11,-30,0,-27,10,14,12,-3,-12,-23,8,0,4,-11,-7,-7,-32,13,37,-7,-30,-11,-14,-14,2,-2,38,-27,3,7,6,-26,8,-1,42,-4,30,-21,-13,-32,-13,29,2,-5,25,-9,5,56,-8,6,-14,1,15,-34,7,-5,8,-18,-4,-5,-6,-10,-15,16,-39,5,2,30,1,17,16,-34,36,-10,15,-15,31,-11,-8,-6,38,-3,-7,-9,-14,5,-24,-24,33,-24,5,-6,13,0,0,33,-32,4,22,10,9,49,11,18,15,15,-6,-36,-46,2,-32,0,9,-21,35,1,-11,0,-3,-11,-7,12,-10,33,-19,0,42,-18),
	(-4,-15,-24,-26,28,21,21,-11,8,6,-24,16,7,-55,-9,-6,14,6,9,-24,-48,23,-9,17,7,27,10,-17,44,5,3,-9,1,37,16,20,-1,-4,5,-12,5,29,-6,3,7,19,0,65,19,2,-20,-17,11,-19,-31,-24,26,-14,-11,4,6,-28,-39,-5,-19,9,0,43,-30,13,18,-35,51,-12,17,-20,11,-32,21,15,23,9,1,-29,-9,-11,-34,-4,26,8,21,34,-19,2,-12,-6,-12,21,26,4,31,46,43,2,-20,34,13,-12,-33,-8,-15,-4,13,-22,11,-1,19,1,0,-30,12,-12,-23,23,0,5,-1,5),
	(0,-4,-4,1,9,19,18,12,-4,-16,-7,-13,15,-40,20,2,22,-24,6,-40,-29,8,10,10,12,11,-37,-2,37,7,-2,-24,13,29,-2,1,-18,-24,-5,-9,5,27,-1,20,13,21,-19,14,2,16,-30,0,31,-8,3,-18,-23,-38,17,-16,4,-19,-37,-16,-19,-6,-4,18,-2,-31,5,-12,-1,-10,10,12,2,1,-2,10,9,0,-4,-34,4,-9,0,-18,33,-7,-10,6,-18,-3,-23,47,9,9,-8,-26,23,-5,48,-26,-24,15,-10,-17,-27,7,-6,-10,26,-18,-8,22,22,12,-8,-5,-15,-8,21,3,-11,14,11,-13),
	(-17,20,-29,9,-20,-8,1,16,3,-3,24,-8,25,-9,-5,21,-25,33,12,-6,-3,28,-1,11,23,-22,-6,16,-3,8,18,13,24,8,-3,12,22,11,4,-20,14,-16,16,-23,3,-13,-8,-10,5,-15,-6,6,10,16,-1,-1,3,14,-2,-15,25,2,-34,-21,-16,0,-5,-20,16,15,-30,28,-18,13,-3,0,18,30,13,-7,6,29,-5,-12,19,-7,-4,29,-6,9,-20,18,-14,-33,14,-11,19,6,11,12,12,-10,7,-2,26,6,-1,22,-18,12,4,-9,0,-28,-7,-24,4,13,1,-9,6,28,17,19,13,-35,39,-10),
	(28,12,19,-6,14,2,-12,-11,-26,-38,-13,16,4,15,16,-3,17,7,-6,22,19,-4,-39,-26,22,-23,-21,-8,36,15,-5,-7,32,-8,-9,-28,17,10,-9,-6,35,26,15,-20,26,-17,2,15,8,17,-4,12,0,20,-21,-10,19,3,6,-18,15,-6,-2,2,-8,15,17,-7,-8,-6,-6,11,38,-4,23,1,2,4,18,-7,-12,6,15,-27,6,25,0,-1,-14,-7,3,17,-18,-30,-2,-6,4,-7,0,-18,10,-3,-17,-24,12,-18,0,-7,-29,20,-15,23,8,-4,-31,5,-4,-8,-23,-4,8,23,-13,17,7,-22,17,5),
	(-16,14,11,6,0,-14,-15,6,-4,-7,19,-9,11,9,-11,13,11,-9,-17,13,-8,2,-8,6,7,8,7,12,-11,10,-14,8,8,2,-1,19,-7,19,12,10,-1,2,9,-13,-15,17,-16,20,-16,2,-4,-19,8,15,12,17,7,14,11,-14,18,-2,-5,-2,17,4,13,6,3,4,-2,-14,3,-12,-14,8,13,14,16,3,-17,-10,-6,-12,-3,-16,16,10,12,0,20,0,-7,-16,18,-9,0,-4,6,6,-5,13,3,-8,17,-5,16,0,-1,-1,-15,-3,-5,17,0,12,9,-7,-11,-5,9,-19,7,9,-9,4,-14,18),
	(-11,-6,15,-3,-17,6,0,-10,-12,5,-17,-1,15,8,5,10,12,7,15,8,-9,-16,16,7,0,-3,-14,5,-9,0,10,-20,-1,11,-19,8,0,0,11,-10,-2,18,8,1,18,6,-11,-7,0,-12,-15,20,-3,-1,-1,-3,14,-10,6,-14,-4,-13,0,-1,19,-7,-17,17,0,-15,16,-2,0,-10,4,0,-15,14,-7,-20,8,2,11,-8,-2,-14,-1,20,-15,-2,6,3,-19,-2,-10,-17,3,4,-16,-20,-2,-11,10,11,0,13,8,0,-6,14,3,-16,-19,15,13,-6,-2,12,-14,-4,-10,17,8,-3,-19,-10,9,-10),
	(-19,-9,-10,8,-3,3,-11,10,13,10,11,5,-6,7,6,3,-19,3,5,2,-13,17,3,-1,-7,-16,3,-1,18,3,-3,17,8,7,7,8,-16,-2,10,6,-4,15,5,16,4,-5,-10,-13,-2,-4,7,-1,-9,-19,13,3,0,9,-10,-4,13,4,-18,3,-7,7,3,-14,8,2,7,8,-13,-5,-9,7,-10,20,16,19,15,-8,-12,0,18,14,-8,18,8,4,-7,21,-18,1,-15,0,0,-8,6,0,-8,-1,5,2,7,5,19,-4,15,-20,20,16,-2,-14,-11,-1,11,-12,-19,-14,-21,-17,3,6,-15,0,0,-11),
	(-35,-8,-14,18,37,-19,-13,-17,8,-8,45,23,7,4,-13,-28,-14,13,5,8,19,-27,-6,9,-5,3,8,7,0,8,0,-27,-23,1,6,15,-35,28,-16,0,9,7,-22,38,-8,47,-4,-9,-42,-22,14,-27,0,24,29,23,-24,0,-8,10,-16,19,12,0,21,-26,-7,-10,3,3,4,12,-37,23,6,-11,-21,3,12,-16,33,-28,28,18,43,-13,-3,-13,-40,34,38,-3,-7,33,7,-8,14,-20,-10,-1,-24,1,-17,15,30,-40,34,-9,15,6,12,3,-5,-1,42,-30,-40,40,11,21,-1,11,-19,18,-1,-43,-6,7),
	(-19,10,-2,9,13,-43,15,4,4,24,-19,0,13,15,4,-35,-29,-28,0,0,5,8,-11,-4,-1,6,-15,-1,14,8,4,0,6,19,-11,36,-1,22,-6,3,-1,2,27,-23,-20,37,6,-18,1,-2,0,-17,28,38,51,-1,-21,7,-8,-2,-2,43,-14,-31,40,-12,41,19,12,3,21,43,-12,12,31,17,-23,28,-33,-7,-6,-1,-23,28,18,-26,-4,43,7,36,-13,37,-5,35,-36,-7,13,16,8,-26,-2,-20,-10,-8,21,-13,-2,-3,17,-29,-24,-1,19,1,5,0,1,20,0,23,11,-21,-2,-29,-40,18,-39,24),
	(-28,14,-3,-8,-5,26,-10,9,-14,31,1,3,19,-6,37,-12,11,-38,-25,-22,-9,-30,3,4,7,7,-13,12,32,4,-17,27,-3,-27,-5,30,-5,-12,13,-19,16,-31,6,-15,-4,29,8,-3,-14,33,15,-17,-17,19,-12,0,-26,-5,2,12,22,-2,-8,-6,-4,-28,35,8,7,-29,12,3,49,35,28,-1,-9,-3,3,-3,1,-8,33,27,15,-7,-22,33,38,15,18,31,-3,1,-21,11,15,12,-6,6,29,0,4,-7,6,-17,-13,33,35,23,-5,-5,21,9,-7,16,33,16,14,-8,-23,3,-24,41,-2,-29,-23,14),
	(-19,-21,-26,7,57,19,-15,16,-1,22,-5,-50,17,-28,24,22,36,-3,35,0,-39,-53,-18,-47,-17,51,0,-9,50,9,5,32,10,-37,-13,24,-39,8,2,-11,-15,-37,39,27,-11,13,25,-21,0,24,-2,-27,-42,-2,-12,-8,-41,18,-9,-20,14,-14,4,-14,-21,-17,23,27,-37,-27,17,15,38,11,35,26,-2,23,6,22,-13,-8,35,-28,19,-11,-26,21,-4,27,2,1,-14,5,-23,46,28,-28,-18,18,10,-32,18,-2,-24,16,0,2,-20,-12,-33,-22,-3,17,-32,19,36,6,-15,7,-32,-16,17,3,10,-15,12,-10),
	(-24,-15,-64,-9,15,48,29,21,16,-7,0,-19,31,-3,42,11,14,0,33,18,-59,-74,-28,-30,-12,51,16,35,48,-6,16,4,6,-42,0,26,-11,6,-2,-2,9,-19,40,7,5,-7,30,5,-36,9,35,-23,-28,-9,0,-15,-32,1,-26,17,-11,19,30,-2,17,-25,22,16,-4,-41,49,35,3,-9,16,33,11,4,-4,0,-25,11,61,-35,-5,-23,-9,24,-19,8,-14,-4,-12,0,-28,17,19,21,-19,-29,19,0,6,28,-32,12,-37,-1,-6,-13,-41,11,-10,-2,-38,33,12,4,-21,8,17,-32,-30,22,43,-14,16,-32),
	(-49,3,-65,-17,28,31,-9,23,-3,-23,-1,-25,-6,-12,22,15,5,17,27,1,-71,-40,-15,-16,-12,2,16,21,3,-7,7,10,12,-29,2,13,0,16,-31,6,-3,-52,21,28,15,-13,33,27,6,-2,-6,18,-7,12,0,2,-37,1,-16,-1,-14,27,10,2,-21,-8,-11,14,-17,-20,30,17,13,11,37,20,-16,23,-11,24,4,3,6,-18,13,-36,1,19,-21,-11,-16,-10,7,-2,-53,-8,-13,-16,-47,5,25,23,19,2,-21,1,-59,11,-26,11,-32,7,28,23,-31,16,22,20,-14,29,16,-17,-27,-28,14,-7,-13,-10),
	(-32,22,-42,18,47,42,-17,16,24,-8,-10,-32,15,-50,31,16,-2,16,5,24,-62,-66,-6,-19,-58,11,10,40,12,-45,-35,10,-4,-36,-14,25,0,29,-14,-3,-12,-59,23,36,-3,-16,34,21,-15,-20,27,-4,-30,-15,-1,-34,-29,-5,-16,-2,0,30,-2,-3,-14,-31,-44,42,-59,-23,48,31,-21,17,10,0,-26,23,-19,25,-5,2,28,-28,44,-44,0,23,-8,0,-39,12,17,5,-31,-13,-1,-2,-35,-11,-13,19,-1,11,-46,24,-23,16,-30,4,-28,-15,8,0,-37,8,31,15,-29,27,-26,-17,-2,3,-16,-43,0,-21),
	(-30,3,-64,33,13,18,-9,42,0,3,5,33,-26,-33,10,23,24,17,33,34,-86,-55,-1,-28,-39,20,1,1,4,-26,-8,-16,27,-27,-2,11,-4,1,-10,9,22,-8,0,8,26,-31,48,14,-3,-9,44,8,-30,-24,11,-53,-9,4,-10,6,-2,30,39,-8,-39,-13,-57,12,-75,-25,31,29,18,12,2,-20,12,39,-23,27,-23,6,17,-52,46,-19,4,20,-2,4,-19,26,46,-6,-29,-37,8,-16,-53,-29,5,0,8,34,-20,22,-42,6,-15,26,-26,-1,34,-18,-40,12,28,16,-38,26,2,-32,-13,18,24,-33,-24,-29),
	(-34,33,-58,-4,1,29,-1,27,15,12,18,20,-7,-61,-5,25,7,-2,-13,12,-52,-25,-9,-39,-21,15,-14,-9,0,-46,-5,-6,9,-9,-18,27,-4,38,9,-11,-1,-3,13,-3,47,-32,25,18,-15,7,11,26,-20,-5,13,-61,-15,-3,-11,-2,2,27,26,-20,-42,-22,-84,33,-81,-45,48,31,0,-4,18,0,-19,20,-28,12,-22,1,47,-42,23,-37,0,25,26,7,-13,26,34,-2,-41,-13,12,25,-24,-14,-3,37,5,42,1,26,-22,6,11,-6,-1,0,27,21,-64,-8,22,3,-9,35,-24,-17,-1,-15,26,-22,-9,-26),
	(-45,14,-52,18,-55,1,21,33,21,0,2,19,-26,-52,4,8,5,15,-20,37,-31,-18,-16,-14,-8,4,10,12,20,-3,24,24,41,7,6,0,-12,48,15,27,4,-20,9,-18,11,-4,13,27,8,-14,9,40,-16,-6,34,-25,19,22,3,12,20,36,25,-27,-49,-2,-27,18,-88,-12,18,16,0,31,-5,11,-10,54,-23,6,-22,10,16,12,50,-24,0,4,-17,5,12,12,33,-18,-1,0,24,10,-30,2,5,13,15,26,-19,39,-35,14,13,-35,-19,4,8,-1,-37,-2,-3,2,0,32,7,-24,-19,-48,-14,-46,-2,-19),
	(-16,24,-70,9,-98,6,0,22,21,23,-3,-15,-17,-63,25,-6,15,41,-3,18,-26,-36,-16,-16,-20,40,17,28,16,-21,39,-1,30,-26,-12,2,-34,16,32,12,0,-4,0,4,39,13,3,0,-11,-12,38,33,22,2,26,-10,11,14,-18,10,6,19,40,-17,-30,-2,-56,2,-98,9,32,44,-8,42,11,-7,-5,31,-15,-4,-6,6,0,-30,44,-11,-7,13,-34,9,28,17,31,-23,9,-10,24,15,-34,7,-5,17,0,37,-1,12,5,17,7,-34,22,-10,19,2,-54,3,1,-4,-4,29,-25,19,11,-55,6,-8,-10,9),
	(-19,16,-64,30,-100,-1,-8,-6,24,21,-12,-48,-19,-50,-2,-16,19,30,-1,24,-25,20,14,-25,-34,7,-4,18,31,-11,1,5,-13,-11,-9,7,-40,12,16,0,14,-7,11,-18,4,18,-5,6,0,7,19,14,26,-9,21,-28,18,7,-13,-16,-1,-11,25,19,13,0,-31,-11,-92,16,19,13,-43,17,0,-25,1,23,-4,-7,-33,0,-7,-62,44,-7,-20,-4,-28,29,35,-19,19,36,-27,-8,45,-29,-16,0,11,3,18,42,-9,14,0,-7,2,-7,-16,-10,19,-12,-65,18,-19,5,-14,-5,-19,28,14,-25,11,-6,-12,-14),
	(-34,-13,-67,34,-112,9,-30,-20,16,16,-3,-13,-9,-48,13,-2,-14,13,-23,-5,-14,-5,21,-22,-34,26,-30,5,-8,-47,-2,13,8,-9,8,16,-33,30,0,-23,16,16,-30,5,14,25,-17,8,-10,0,5,12,11,-22,23,-45,33,0,9,0,16,-5,9,5,-28,-19,-27,19,-86,25,28,19,-34,14,-4,-10,-1,38,2,-1,-32,3,18,-53,17,-15,-9,0,-17,-8,35,18,33,22,-21,19,5,-37,4,-22,16,2,-19,21,14,0,-2,-12,-53,-5,-13,12,1,-13,-45,14,17,0,-19,-9,-9,0,26,-42,-29,19,-5,8),
	(-32,1,-50,31,-39,9,-4,-4,29,11,-31,-18,-40,-31,-24,-17,0,33,7,25,-27,-15,18,-20,-20,6,0,-4,-17,-4,14,4,16,45,-2,36,3,33,-24,15,31,5,-37,0,0,23,-33,32,4,-25,10,0,2,-30,16,-19,25,17,-14,-18,4,16,44,-10,-33,-17,1,19,-46,34,20,23,-33,-18,33,-27,-7,7,-43,1,-5,6,-21,-44,40,7,18,1,-1,-12,19,14,34,36,-5,16,30,-9,0,5,8,8,-12,19,-21,30,-3,-44,-48,-14,-11,27,21,8,-31,50,-3,4,0,15,-2,4,-2,-21,-49,2,-27,18),
	(-29,19,-8,54,-12,12,17,7,25,34,-4,-17,-28,-15,-34,-7,8,15,-5,4,-38,-13,14,-8,-16,5,-3,0,6,-20,-5,-10,4,18,19,43,-5,46,-25,-5,1,28,-40,-20,16,29,-33,8,9,1,-2,32,-12,-27,5,-43,18,-14,-11,-16,-3,21,19,7,-27,-8,-27,14,-61,-17,20,27,-51,-36,16,-31,-7,30,-26,-6,-28,6,-4,-39,50,-36,8,-10,15,-10,7,24,28,7,-25,30,11,-20,-2,20,6,20,24,49,-9,19,-13,-28,1,-13,2,15,30,0,-6,37,6,-5,2,-9,-18,-25,-30,-30,-15,37,-18,1),
	(5,5,-2,15,22,16,20,-31,7,30,4,-31,-29,-38,-52,12,2,46,17,31,-39,-19,9,-12,3,33,-47,-10,-11,-32,7,1,40,8,28,30,15,26,2,15,14,26,-74,-20,8,5,-33,14,-8,8,-7,42,-19,-6,-17,-38,3,18,14,-16,21,15,34,12,-1,25,-14,35,-17,-8,10,0,-12,-58,12,4,19,1,-30,-8,-23,16,0,-47,13,-6,-3,11,8,2,6,25,-17,31,1,4,-31,23,4,-5,-2,2,22,46,-23,13,13,12,-39,10,4,0,15,-2,26,50,7,-8,-6,-22,22,-25,-25,-31,-22,35,20,-11),
	(-7,19,-22,24,9,-7,10,-47,21,23,-16,-26,-33,-17,-37,6,7,26,-6,36,-18,-18,16,-25,-10,13,-11,-31,-1,5,21,-7,17,30,13,-4,-11,5,0,25,13,-4,-69,-16,20,-2,-41,19,-6,-11,-27,33,10,18,-6,-43,-10,-16,1,-18,1,48,-4,-20,0,9,-8,21,-16,2,-1,21,12,-63,-4,-12,4,31,-41,6,-11,25,-4,-13,41,-4,18,27,-6,-13,10,6,-14,-1,-46,34,-23,15,-1,13,33,-13,40,27,-11,23,-1,-11,-6,-1,-4,19,16,-2,41,7,23,18,-14,9,14,3,-37,-17,-9,21,0,14),
	(-27,7,-5,7,65,0,-29,-20,-3,-12,3,-6,1,-23,-15,32,13,2,18,20,-17,20,24,2,0,2,14,-37,-4,-13,-7,-24,-18,17,-5,34,-17,9,-18,15,-10,31,-28,-11,25,-12,-15,6,26,2,-2,11,-21,7,-9,6,-23,-21,-13,-14,10,13,11,25,11,21,-10,9,-27,20,6,-1,-29,-85,32,-1,-7,-4,-31,6,12,15,-13,19,4,2,0,27,6,-28,0,-8,-7,-25,-58,3,-63,5,20,21,21,35,34,24,-6,-1,-6,15,-6,-5,-4,0,3,-13,3,-7,23,-23,-38,4,-3,-20,-25,18,7,33,11,8),
	(7,38,-12,6,38,7,-2,-20,-5,13,15,-17,-20,-27,-31,-5,14,0,4,-5,-54,7,33,-9,-16,-1,32,-8,17,0,-11,-5,-4,27,11,14,-10,-5,-26,-1,-10,2,-20,0,30,-24,-1,-4,-2,-15,0,12,-2,10,-2,1,-24,-13,21,4,3,25,-9,5,-49,-8,-3,16,-9,21,-7,-21,-18,-63,0,-23,2,-23,-22,-2,-1,-1,8,-7,9,-11,19,22,0,-29,-22,7,-19,-11,-6,-12,-61,6,2,24,23,14,22,22,-13,0,-14,-33,-2,11,7,19,16,-10,13,-1,14,-29,-16,-4,22,-15,-52,15,0,32,28,-5),
	(-10,42,-4,-35,38,17,-9,15,-51,-25,-23,-17,-22,-3,-16,0,13,-12,40,6,-27,-8,0,-12,13,-1,4,-38,-13,9,-15,-19,-13,16,7,0,-7,6,14,3,0,11,-10,-18,23,9,13,30,52,21,-42,-15,-30,-11,-20,-7,10,-13,-1,8,-10,-6,-12,0,-72,34,23,7,2,14,-20,-1,-13,-19,34,-38,-4,-19,2,-11,28,-6,-22,20,-23,-16,33,7,14,-16,14,0,5,-33,-4,0,-29,-3,32,30,-4,20,-10,5,-11,-17,-14,-39,-14,5,-19,4,15,21,23,-41,-4,6,-43,-9,15,11,-52,-4,-15,31,-14,11),
	(-7,35,19,-20,38,10,-25,21,-6,-3,-4,1,8,-33,-8,-9,21,-27,38,-18,-21,23,34,12,15,-21,10,-9,19,-20,8,-5,20,17,8,-7,-5,-14,17,-1,41,8,-34,-18,3,22,-21,-27,21,25,-8,-2,-9,18,2,2,16,-1,13,-7,-9,-14,-30,9,-98,23,12,-6,24,23,-26,-21,-18,-31,8,-42,5,-5,17,10,39,11,15,15,11,10,-1,-11,0,-7,-3,15,-2,-12,17,22,-37,5,-5,33,6,-1,7,-3,-31,10,1,-50,-6,35,4,11,6,17,28,-32,5,25,-20,13,2,-18,-59,-5,11,7,11,-27),
	(30,-6,-2,-46,16,9,-1,34,-47,-34,-1,25,-1,-4,-24,-45,-21,-11,25,-56,-17,27,3,-8,12,12,3,-20,-6,-2,0,-31,5,26,41,-12,26,-2,31,0,31,22,-9,-18,11,6,-21,38,31,8,-15,-13,0,-1,-22,-2,8,-50,3,-13,-20,-27,-54,6,-66,22,22,0,22,-2,-29,-33,32,-19,7,-35,23,-9,11,-2,60,7,0,-1,-36,4,3,16,23,-29,8,8,-30,-25,23,4,-1,-3,9,17,23,27,17,-15,-13,-9,22,-24,2,27,-29,0,18,-18,50,-22,-19,18,5,-25,19,44,-46,9,9,-34,7,-24),
	(-11,-57,19,-33,-55,6,-15,23,-9,-66,-35,35,31,-18,1,-40,-10,-6,10,0,-44,6,-42,-12,27,6,-11,-23,15,-11,16,-21,22,-22,27,6,30,-4,20,20,40,44,-5,-45,66,-3,-26,41,40,8,-11,18,11,11,8,-2,35,-21,-1,-7,4,-33,-54,-1,-31,53,24,-11,39,23,-3,-1,18,-16,-4,-15,67,0,26,-2,21,38,-24,-28,-30,-13,32,-9,9,6,-27,-13,-10,-33,33,29,4,-15,-4,-7,5,57,-23,6,19,7,22,-3,-6,-13,9,-18,22,-1,46,-36,-5,29,-21,3,25,5,-32,-20,-16,-55,-12,23),
	(0,-28,-11,-1,-32,4,-15,37,-5,-58,10,58,9,-4,5,-14,-8,5,44,13,-10,27,-49,22,30,20,3,1,-6,-15,12,-34,41,-1,43,5,17,25,-18,-4,15,19,24,-35,70,-2,2,31,25,0,-30,14,1,36,5,22,43,-45,13,-8,7,-19,-28,-40,-46,32,21,-25,37,3,-19,-14,-27,-22,-31,-10,65,-8,4,20,-16,44,6,-11,-7,-38,14,3,2,1,7,7,12,-42,32,30,10,-10,-18,37,-4,48,-28,19,32,8,18,1,-4,15,6,1,8,2,44,-23,2,47,2,5,16,-5,-12,-13,-48,-7,3,-3),
	(33,-5,0,-8,-17,-14,4,8,9,-24,-6,53,14,-44,-2,-10,-21,30,30,13,7,-11,-10,9,45,-4,-31,10,-16,-7,15,-12,1,4,-4,14,-13,-17,-9,-30,20,29,44,-16,38,-11,7,14,17,25,-19,2,32,28,0,-1,48,25,16,10,35,-18,-16,-3,-13,27,0,11,-8,-19,22,-14,27,-6,11,-11,44,20,-26,16,-34,32,-42,-24,6,-44,43,-8,-7,-25,-15,28,-18,-48,36,14,-16,0,-5,18,32,52,39,14,14,-3,10,12,-22,1,22,8,27,40,2,17,18,37,-30,3,52,-14,21,-6,-21,0,12,8),
	(40,12,-15,-16,6,23,6,-15,-11,0,-13,6,-16,-34,12,22,-1,-14,-7,-26,0,-3,-4,-21,1,17,-8,16,18,9,-33,4,2,-3,-4,-6,-8,-4,-10,-5,-17,-1,5,13,18,8,40,-13,-7,28,-35,-25,-7,1,4,-21,-19,8,-1,-18,-15,-7,-19,-4,-3,15,-2,33,7,-1,17,-23,14,-9,7,7,8,-9,13,19,9,4,-3,-28,-24,-21,-11,4,13,7,10,26,-6,-10,3,13,2,-10,26,34,6,46,8,-28,-17,10,-4,0,0,13,10,-2,21,3,-45,37,16,2,0,-6,16,-25,-8,-9,12,18,26,13),
	(-15,13,-17,-17,-20,0,15,-7,-3,13,-20,-19,-10,4,-7,-12,0,-8,-11,7,-20,18,9,16,-11,5,11,-5,14,-17,-14,-1,-7,11,-15,19,20,11,-3,-3,-17,1,-19,11,9,-8,8,-5,0,11,-19,1,-7,-20,0,-3,5,0,8,-8,-10,6,-16,-13,2,-16,6,-8,-19,-16,16,-12,10,-9,-7,-10,-6,-12,18,16,13,1,-13,0,-15,-9,13,0,10,17,10,0,-10,17,-13,1,-15,0,12,0,14,-19,17,12,-2,-16,-18,-7,4,13,15,-5,0,2,-19,0,-5,0,-1,10,11,15,13,-17,-4,3,-14,4),
	(16,-4,12,-1,-17,10,-20,-15,-13,-5,18,-1,4,-8,3,5,5,8,-17,-17,19,-16,0,8,0,6,-10,-2,-8,-4,5,16,-16,-19,1,4,13,-12,8,-4,-18,-15,18,-13,17,-2,14,-17,8,-12,-11,-13,11,17,-3,20,3,9,-2,14,-6,18,-13,-14,11,-18,-8,2,0,-18,-14,-17,6,-5,-5,-8,0,20,-9,0,4,10,8,8,-15,17,6,0,-10,-1,-13,-6,1,-19,-14,0,12,-14,-7,-20,5,-10,0,5,-2,17,13,16,-15,19,-10,-5,-7,-8,-15,-5,13,0,-19,18,-7,7,20,4,-2,-13,6,-11),
	(-9,-17,-20,46,4,18,-8,3,40,2,16,5,36,36,0,1,-16,5,13,2,0,-28,14,23,0,7,13,17,19,-3,1,14,-24,-14,-17,45,-14,-1,6,-11,-22,5,-24,11,-34,11,15,17,-28,-15,-14,-23,-3,-10,22,-21,-11,-9,-41,-16,5,22,29,26,52,-7,6,-16,1,15,32,23,-4,-5,13,-12,-14,-8,6,-40,19,-10,-6,34,36,6,9,-2,-31,31,0,-9,-8,38,-42,-36,-8,0,2,-29,-14,4,-5,32,24,25,8,-56,-9,-6,0,4,-25,12,9,1,-21,24,30,4,-20,10,2,14,-16,-17,-3,8),
	(10,-8,-20,-4,-28,8,7,3,8,-20,15,-18,16,3,-8,-4,1,27,13,4,-12,-8,7,31,2,9,0,-10,17,8,32,-15,7,-8,-27,-7,-7,9,-6,-10,-13,-8,-3,-11,-4,4,-20,26,-8,-35,-15,18,-3,-2,40,31,-32,12,-14,13,-12,14,-11,-9,0,-21,30,-32,-20,7,8,17,26,23,-5,15,9,4,-16,23,0,3,-9,9,-4,-50,-37,22,-2,5,-24,16,-22,17,-15,5,11,13,6,-26,17,-19,7,26,6,3,-20,-46,0,15,-13,-7,-8,-12,17,-14,3,8,1,-15,9,-3,-25,-6,-6,-30,-10,-6),
	(-42,10,-25,-24,-11,40,24,-28,-4,29,11,-30,45,-15,42,9,17,-17,7,18,-64,-70,8,-23,-21,29,-46,-17,33,-26,4,28,17,-50,-23,8,6,-32,-6,-26,-21,-47,61,32,0,5,30,-1,-20,-5,12,4,14,-20,26,-13,-36,0,-8,-11,32,17,-10,14,-7,-39,53,6,-13,0,10,5,46,34,26,17,-36,22,-5,13,2,-31,38,1,1,-23,-43,8,-6,43,-45,-15,-23,-29,-16,11,45,5,-44,37,1,-22,7,34,12,6,-10,30,-13,-5,-19,5,10,-18,-44,-12,41,-21,-3,13,-11,-36,-18,32,39,-28,-2,-3),
	(-23,2,-34,-14,60,18,-15,-25,24,15,-20,-22,43,-26,40,-31,-12,-4,71,13,-32,-87,16,18,-39,-30,-9,-24,39,-5,-21,32,-25,-38,-23,-5,-4,16,-6,3,42,-24,11,16,-28,9,49,-5,-4,32,-6,-5,7,19,33,19,-24,21,1,-5,-1,4,-8,-2,-44,-36,20,-34,-27,-19,3,39,51,3,50,-9,-52,-7,8,4,-28,-56,13,36,-7,-10,-5,23,-9,36,-39,-4,-19,-17,-36,11,49,-11,-19,16,12,-49,-22,9,4,-35,4,13,-9,14,-32,-9,-13,8,-31,-34,-21,19,-33,14,0,-16,1,13,23,-53,-20,22),
	(-56,5,-26,-6,55,16,10,4,19,21,-5,1,6,-56,26,-16,5,0,25,15,-72,-41,0,24,-23,-17,34,-34,32,-26,-13,-1,-23,-64,-24,17,-2,10,-18,2,40,-18,11,1,-43,22,15,3,-10,9,5,3,4,-2,24,7,-10,3,10,-9,-12,10,-1,5,-44,-21,13,-21,-19,-30,21,25,29,-4,35,-18,-22,-1,14,-3,-6,-49,37,2,3,0,-22,3,-27,44,-43,-9,-12,-11,-19,-12,31,-20,-43,7,24,-6,-7,6,-36,-16,7,20,-1,9,-19,-23,-31,25,-3,-18,7,36,-4,23,-6,-42,4,-6,43,-56,0,-4),
	(-37,-5,-21,-19,68,-11,-2,44,18,18,3,5,10,-17,28,9,-13,11,56,13,-30,-64,-33,-12,-40,8,34,-7,41,-25,-47,0,6,-76,-26,23,-6,10,-7,9,-6,-36,4,0,-20,24,19,-29,12,-2,37,-19,7,14,-3,-22,4,16,10,-15,-5,0,-8,11,-32,-27,14,4,1,-24,4,43,17,11,8,-27,-3,-18,17,7,-13,-14,21,21,18,-42,0,-16,12,26,-53,6,-1,-47,-43,3,20,14,-31,25,-12,-16,8,3,-15,-31,-33,28,23,3,-19,-23,11,10,10,1,20,8,-12,2,7,-41,-5,-17,11,-21,-3,-16),
	(-57,13,-33,-2,55,-21,3,-1,0,10,-12,4,-26,-34,59,2,3,-1,21,5,-57,-46,-14,-39,-38,-13,-7,0,2,-57,-36,-20,1,-21,-9,0,37,-12,14,-11,-7,-14,28,8,-12,0,24,-26,-1,-1,28,6,0,-9,19,-15,-29,26,19,14,-3,7,-13,-5,-45,0,-13,1,-39,-35,-16,14,-7,6,-7,-32,15,-12,25,33,-21,-27,-9,-5,3,-10,0,-7,-1,15,-49,-19,24,-31,-8,-32,-6,27,-40,9,-9,23,3,-13,8,-27,-28,35,-3,7,-11,10,-6,21,-28,-19,-10,8,-13,5,11,-4,2,19,30,-24,-3,-28),
	(-60,-10,-12,-32,47,-7,2,2,18,16,-3,22,-6,-31,33,-12,-5,1,0,25,-38,-33,15,-38,-39,4,21,-7,-17,-7,-11,6,-16,6,15,-15,3,-9,-7,25,11,5,5,-29,3,-6,7,12,32,13,16,22,-6,-23,16,-25,-6,4,28,10,3,11,5,-13,-79,13,-17,-24,-40,-37,-14,4,-15,17,-4,5,9,-10,22,30,-17,9,21,17,0,-17,30,5,-7,11,-29,3,27,-41,13,-20,24,42,-69,33,-30,4,-16,-7,-8,-6,-7,1,13,2,4,-6,-2,-10,-41,-11,9,1,-15,31,10,2,18,-1,16,-4,19,-29),
	(-33,10,-50,-12,9,-27,-26,33,-18,-11,11,18,-41,-13,-2,27,-14,22,-10,-4,-49,-14,24,-34,-4,0,15,0,-14,2,-10,-4,19,-2,-5,4,10,-7,-8,2,-7,-8,-10,-7,3,4,8,9,7,-11,-12,-6,4,-25,21,-16,-18,20,4,10,-2,41,10,-39,-54,-15,-49,4,-37,-12,-3,4,17,-9,-6,-18,14,17,16,0,-2,38,3,5,27,-23,-1,24,12,19,2,14,55,-10,-3,1,14,11,-28,12,-8,20,1,-10,-1,-31,8,-14,0,-25,11,1,4,-10,-29,-35,-11,-13,-2,40,0,-2,-7,7,-9,-24,5,-28),
	(-25,7,-38,-12,-96,-10,-16,17,28,-6,-11,22,-42,-60,-11,24,0,29,0,-5,-46,-40,9,-1,0,6,9,-8,-21,9,-4,18,36,-3,-11,0,-13,0,22,-18,5,-12,16,-23,34,-9,8,-7,9,0,-10,28,5,-15,32,-10,23,15,19,-7,15,31,1,1,-33,-5,-33,-11,-67,4,-8,-16,-1,6,-8,18,35,19,26,7,1,30,-26,3,18,-14,18,7,26,-5,2,26,29,-27,44,22,53,32,-15,13,-13,1,-12,2,-1,-4,23,-14,26,-31,11,36,0,-7,-16,-28,7,2,22,35,14,24,4,-18,-9,0,27,-10),
	(-53,-12,-22,6,-97,-9,10,26,19,2,-20,-10,-7,-44,-8,-10,7,10,-6,0,-38,-34,-20,-6,-29,29,13,20,30,-20,20,7,20,-8,7,5,-10,33,37,-21,-5,-14,14,-23,29,0,-7,31,0,17,23,24,15,-2,1,-20,17,5,27,2,8,30,-8,-6,-12,12,-48,17,-43,0,8,-16,-14,27,24,3,-2,31,36,9,3,26,-29,-29,1,-10,-1,-13,-2,3,17,7,33,-11,18,8,57,21,23,0,-12,3,-28,25,16,1,34,-26,-14,-8,9,15,-3,4,7,-35,5,-8,18,-8,1,22,-5,-14,-10,4,-3,-6),
	(-47,12,-60,7,-108,-22,25,-20,40,0,13,-13,-4,-46,8,12,-13,29,6,23,-25,0,-17,1,10,-5,-64,9,17,-2,-3,-4,34,2,5,3,-1,19,18,0,20,-9,-3,1,21,15,4,11,15,15,-12,-13,29,0,21,-13,17,19,10,-10,-15,7,27,-17,-16,23,-5,5,-39,0,-14,10,-53,9,-1,6,13,25,-6,4,-23,20,0,-63,28,-40,13,-5,1,6,13,2,39,5,15,28,43,5,10,-7,0,-7,-7,35,4,10,26,-4,-13,0,-10,14,12,19,-33,1,0,0,9,16,1,28,-4,-13,-42,8,-8,-6),
	(-33,10,-53,25,-38,-6,-12,-16,30,5,-14,6,-2,3,-9,0,-21,30,11,-8,-62,-6,9,-15,6,-10,-57,31,-10,-4,0,-24,16,12,15,-7,-12,32,21,-22,-2,23,-30,1,25,41,-9,18,30,-11,-4,5,22,-10,1,-10,-12,20,-17,1,-16,21,26,9,-11,6,-18,9,-47,6,-5,-9,-31,17,-2,-19,0,39,14,13,9,24,-30,-51,-3,2,-8,-13,-11,0,31,30,27,23,1,-8,19,-5,36,-8,-8,-16,-32,26,12,26,11,-23,-8,9,-14,9,13,24,-1,10,1,23,7,9,6,7,-6,-30,-31,24,-18,-10),
	(-19,2,-51,29,4,-17,-10,-5,42,10,-18,-34,-20,-25,-10,-20,-10,22,9,21,-57,-9,-15,16,-16,18,-43,18,0,0,10,-7,0,7,-19,16,-5,19,-8,-26,11,12,-3,-9,9,40,-3,-4,4,3,-1,19,5,-24,5,7,18,25,12,-21,-21,18,15,19,1,16,-17,-21,-22,-25,21,0,-19,1,-5,8,9,24,-15,5,-12,-4,-8,-29,22,-7,-29,-4,2,20,32,-6,20,20,-16,15,20,-22,37,3,6,-49,-13,0,-20,20,6,-6,-7,20,-6,-14,25,-6,-20,27,-15,-2,-14,2,7,-12,5,-21,7,30,-7,-5),
	(1,-1,-44,28,43,-5,0,-19,11,-15,-4,0,0,-16,-20,20,-19,23,18,12,-42,-31,-23,3,0,12,-48,1,10,7,15,-28,20,-5,-6,26,-23,36,-42,9,5,31,-53,-21,14,19,5,-12,22,-2,-18,16,-5,-41,16,14,-18,28,-22,-11,-24,10,28,-8,-29,-6,-16,2,0,-32,7,16,0,-16,4,-7,0,32,-21,7,-45,22,0,-18,0,-20,-11,25,-12,3,22,13,11,24,-30,-14,27,-3,14,-4,-1,-34,15,18,-7,27,-1,8,-16,-25,-21,24,31,22,18,41,-9,10,0,19,21,-16,4,-12,-14,31,-10,1),
	(9,7,-29,25,57,20,6,-5,10,-17,-8,-3,7,-45,-16,8,10,34,-7,-16,-68,-14,4,19,-9,11,-6,8,-15,9,3,-8,36,25,-9,18,-22,13,-14,-3,18,9,-70,-37,39,-27,11,-7,21,-12,-21,13,21,-35,12,8,-14,-3,-12,-6,0,0,34,-1,-11,28,10,-3,3,-19,-17,0,-42,-50,6,-22,16,20,-8,18,-29,-2,10,-7,11,-26,27,0,2,-24,-22,5,-11,-6,-28,6,-8,-11,-13,-26,24,-11,14,1,-9,-1,-12,-27,0,8,12,-3,29,0,-13,40,13,5,0,2,6,11,3,14,-40,29,-4,-4),
	(21,0,-25,37,37,-3,0,-16,-11,25,21,-13,22,-22,-45,1,36,37,17,28,-65,3,32,8,-8,3,5,-5,-12,2,20,-24,39,29,3,-8,-22,-18,-33,-1,9,19,-62,1,0,-22,-27,-19,19,13,-25,16,-16,8,7,-2,-18,1,23,11,-7,8,40,12,-10,-5,-14,29,-5,-37,23,-8,-28,-40,25,-15,20,36,0,0,-7,-11,9,-16,39,20,29,0,-16,0,-5,26,-11,14,-20,14,-29,5,13,-13,5,-5,49,3,-11,20,-1,-19,-5,3,-22,14,-7,19,1,27,24,-12,-17,12,11,-6,-12,14,-13,44,29,-7),
	(35,9,-39,32,48,3,-11,-12,-11,-3,8,-16,29,-55,-39,0,29,2,17,20,-57,-12,61,0,11,11,23,-7,25,2,15,-23,11,21,-15,39,-18,14,-48,-8,4,2,-50,-17,6,-8,10,-15,17,12,-5,-2,-22,-7,6,3,-4,9,-1,9,21,8,-3,33,-16,-10,-12,24,-3,-22,29,-13,-34,-53,25,16,11,-12,-1,-17,-13,-23,5,-8,21,-28,-5,-5,18,-40,-31,35,-30,-21,-62,-10,-19,-16,6,-2,13,0,56,15,-5,11,-14,-20,-11,-14,-17,22,31,12,4,17,14,1,-31,-13,-1,0,-29,8,-37,42,-6,2),
	(28,-9,-8,-2,30,30,2,-6,-2,1,-19,-28,8,-15,-26,35,28,23,23,-16,-33,-23,26,-5,16,31,-3,-29,19,9,23,-11,19,36,-4,23,-16,2,-21,5,3,35,-21,-1,30,-41,-29,-4,15,-13,7,21,-44,-11,-19,-2,2,-12,-12,4,0,18,-9,-5,-29,13,0,24,15,7,3,-7,-6,-72,4,-17,16,19,-22,-18,34,23,-4,-12,39,-23,1,29,13,-69,-31,22,-69,-22,-47,5,-62,16,-6,-8,-7,21,38,49,15,5,0,-45,-26,-15,8,21,33,0,12,18,18,-1,-28,9,11,-14,-44,13,-20,1,17,-21),
	(-9,22,-8,13,27,25,-20,22,-40,0,20,-1,10,-9,-41,31,12,33,23,-12,-39,24,22,-9,-6,-4,41,-19,-23,-2,21,-36,-4,27,2,23,0,7,-13,-11,-2,2,0,-8,21,-21,-24,-16,6,9,18,24,-20,5,-3,20,-13,-14,-34,5,10,-5,-1,15,-60,-12,-4,27,3,-4,8,25,-15,-58,27,-39,16,17,-16,6,-6,-27,-13,-3,32,-33,-14,-15,4,-34,-14,5,-72,-40,-25,-6,-61,-13,-5,28,-18,16,-2,43,5,37,-4,-54,-13,10,-18,7,36,-32,27,7,-18,16,-24,-10,17,-1,-54,3,-32,-3,5,1),
	(11,-1,17,-18,17,-7,-49,16,-49,12,23,21,0,-8,-36,38,28,8,-2,-5,-30,11,43,5,4,1,39,-11,-28,21,15,-11,-14,-9,8,1,-17,-2,-12,15,0,16,-23,-16,19,-23,-16,-23,15,14,42,4,-22,4,7,4,-3,13,-27,-2,-8,22,-20,8,-70,2,-12,1,0,-26,0,3,-27,-34,2,-17,-13,25,-26,-5,17,-12,-15,20,29,-15,27,9,-21,-8,-13,-19,-58,0,-21,-14,-71,-24,-9,1,-6,24,30,22,-25,25,-25,-41,0,2,-30,37,13,-29,38,-17,-3,4,-6,4,16,5,-25,-14,-19,-14,17,-11),
	(24,-30,4,-33,12,36,-50,33,-23,6,17,50,2,-30,-31,14,35,-3,-1,-33,-64,-4,14,-36,-19,-20,25,3,11,17,-19,-2,-6,-1,6,7,10,2,5,-11,30,39,-8,-11,26,22,-14,-4,9,23,-20,-12,-42,-5,-14,-15,-3,0,-28,4,-21,17,-32,-6,-22,3,0,7,43,19,-13,4,2,-19,0,8,8,-24,4,15,35,-14,4,-1,-20,0,16,8,14,-24,-4,-5,-81,-28,-8,-29,-42,-11,23,44,4,15,16,12,-43,10,-34,-62,0,11,-46,38,25,-26,18,6,12,13,-20,8,32,14,-24,12,2,-24,1,8),
	(17,-68,0,-24,6,30,-30,12,-2,-32,-18,56,9,-28,-13,-17,13,-1,10,-36,-61,22,-16,-26,7,11,11,-27,-15,8,4,-18,-22,21,16,0,22,0,-5,-25,27,29,-3,-15,17,17,-16,8,5,22,-45,-9,-36,22,-10,6,21,-2,-35,-17,-34,-38,-90,13,-34,30,-27,27,41,-12,0,4,-10,-33,13,-20,-2,-10,-10,-17,32,-11,3,19,-12,-19,46,15,-10,4,-4,-3,-31,-45,11,3,11,-34,18,0,19,48,-11,19,-36,-13,-18,-35,-18,23,-36,-3,18,-9,17,3,-10,-3,-31,-25,39,31,-15,-15,5,-37,-13,4),
	(19,-29,-3,3,-37,8,-10,24,5,-66,-6,55,28,-36,-1,14,-12,-6,21,-5,-35,-18,-18,-12,8,13,0,-4,-3,22,11,-23,21,0,23,42,27,25,-22,-6,53,12,15,-13,43,3,28,35,19,15,-30,36,26,56,27,18,24,-5,-7,-21,11,-10,-54,-11,-32,45,-5,-6,-1,7,2,8,-27,-16,4,-29,59,0,7,28,4,32,-14,-47,-26,-18,53,-4,-29,-36,-12,44,-33,-41,17,-4,-10,0,-10,43,24,57,15,0,-11,24,13,-2,-20,-4,-5,-23,47,12,7,-41,27,65,14,38,37,16,-6,-15,-28,-22,33,-14),
	(36,-1,-3,-36,1,-3,0,20,-5,-19,-11,39,-2,-6,-35,13,-24,-1,10,-40,-23,-2,-27,0,-2,11,-7,-20,32,34,-15,-20,24,18,-10,-11,22,-6,-29,0,35,59,27,4,25,-26,43,14,6,10,-37,-16,0,1,-24,0,38,-30,-17,-6,34,-37,-35,-4,-19,38,-14,36,-12,12,-9,0,31,-6,27,5,34,0,8,1,-1,39,-16,-44,-21,-29,25,-9,-33,-27,-20,15,3,-40,12,1,-25,7,32,14,25,54,1,-17,-8,20,8,13,-42,-21,3,-30,14,18,-15,18,44,30,-18,44,3,-17,-8,-1,-17,20,24,-9),
	(25,-14,11,-12,16,31,33,3,-16,-3,-7,10,-12,-34,0,-14,8,-38,-18,-39,-36,-15,-7,-9,-19,9,-19,-14,19,34,-22,-17,1,19,-32,14,20,-9,-3,20,22,-1,29,9,38,1,30,-1,-6,31,-31,-11,-3,19,-29,-29,18,-26,-19,-15,-24,-18,-23,13,-15,21,1,25,-10,0,3,-30,21,0,-9,16,25,-6,17,-7,3,-1,2,-8,-18,-23,17,12,22,-17,-8,2,-9,-7,16,-27,-3,4,1,27,41,40,19,-35,-35,-11,9,22,-3,29,-24,-17,14,3,-33,0,4,6,-14,9,23,1,21,16,10,4,32,-7),
	(-14,7,-13,-10,-12,5,3,0,-12,17,-10,-10,-13,-7,6,11,14,-8,8,8,-10,9,-2,7,-18,-13,-1,-14,20,14,8,-5,15,-7,-18,20,15,-17,18,6,0,-5,-1,-8,2,18,-13,3,-11,-1,10,10,-1,-5,13,14,-4,-14,-14,20,-13,-15,4,-19,-17,7,-6,16,1,18,-1,3,-16,-7,0,19,17,1,8,-13,0,12,-9,-1,-20,0,-18,-11,-1,-18,16,10,-7,-17,0,-9,14,-15,19,-11,20,-13,18,0,-16,15,-13,6,0,14,-7,8,14,20,-14,-18,-17,8,-11,-2,12,-8,-15,1,-20,0,6,13),
	(2,12,2,-6,-4,-4,5,-2,12,4,0,-12,3,-21,-5,-3,4,10,21,-3,-29,20,16,-7,-32,4,-8,5,34,33,-13,15,10,0,2,29,-24,16,8,19,29,9,-9,0,-4,7,30,-14,2,11,18,2,-5,-27,29,-9,7,20,-15,-6,15,33,-3,-9,0,4,-8,18,4,-17,-4,2,24,5,30,-1,-24,3,-15,-1,1,-1,-10,25,31,-1,-11,31,-2,3,16,2,-1,-8,-27,1,-5,0,0,27,-8,8,0,12,11,12,-25,7,18,-19,-30,7,22,20,13,7,-6,1,-22,14,3,10,-6,-20,6,-21,-18,9),
	(10,-17,27,-7,-15,-46,-6,6,8,22,-17,31,7,2,-12,-12,8,-16,2,12,7,2,-31,-9,13,-10,2,-2,-1,17,-30,-16,21,-31,-6,7,12,-9,17,38,14,0,7,-18,-6,21,-1,-17,19,33,13,14,18,-3,7,4,-17,-5,30,-1,-20,8,7,-14,-19,32,19,22,28,16,5,5,19,31,-4,-12,-23,7,15,14,-21,-13,4,50,-1,3,33,8,20,9,-2,-14,39,-19,6,-20,33,10,3,41,2,0,7,6,9,-43,-14,23,0,25,-20,-20,-3,33,31,-5,-23,12,-16,14,29,-12,-16,26,0,17,-18,0),
	(0,1,-11,-26,-2,-9,-11,6,13,15,22,-23,34,25,-2,-25,21,3,33,28,27,42,0,30,-1,-9,-28,-23,30,20,-4,-3,8,-37,-20,10,15,-5,-22,7,-19,-40,0,0,6,1,25,-15,-18,-10,25,-31,-10,-6,25,17,-10,15,16,-14,10,34,17,9,-40,0,10,-3,0,-4,3,3,40,16,5,31,-4,13,16,25,-12,-19,40,21,1,1,-10,10,-5,-5,-28,-8,-14,7,15,-12,47,20,-13,7,0,-30,-3,-24,3,-21,-33,15,4,0,6,-12,-13,0,-6,-24,3,24,-25,-2,6,-10,-38,38,17,-17,-11,-22),
	(-24,24,-21,-31,-16,42,25,9,5,13,31,-21,6,-1,13,-19,33,8,13,16,0,28,10,4,10,0,-11,10,38,4,-24,-10,17,-48,-2,-16,-3,-5,12,26,1,-49,2,-9,6,-6,40,-35,-17,3,2,1,-12,13,7,-4,-28,25,-21,19,-10,-4,4,4,-32,0,36,-13,-1,-13,-9,-5,47,-10,32,14,-24,-6,1,23,-4,-39,44,-3,0,4,20,25,15,15,-24,0,5,-25,2,-1,34,33,-48,-2,18,-29,-22,-17,-18,-17,-24,44,-15,-11,-3,-18,11,25,-41,-10,5,26,-24,29,-7,2,-26,22,36,-36,0,-6),
	(-49,11,7,-14,65,8,-4,0,-8,18,8,17,8,-29,14,-7,-1,7,52,4,-27,25,0,1,-5,-13,39,-14,13,-32,-44,-6,14,-28,-12,-16,42,15,11,16,44,-56,8,-15,1,0,22,-56,42,21,16,19,-7,-12,0,11,-21,-5,8,6,12,25,17,-32,-19,-2,43,-37,1,2,-47,10,13,-7,0,22,-31,-14,6,0,-7,-42,32,-27,6,-2,39,26,1,18,-10,-17,3,-22,-37,-11,26,8,-25,5,-26,-27,-33,-22,22,-22,0,10,6,31,-32,-6,-13,40,-19,-21,-3,11,-27,31,23,-1,-36,45,41,-22,4,-12),
	(-42,8,-35,-20,60,-35,10,2,28,30,-31,10,20,-9,39,-8,-20,25,40,24,-4,-27,7,14,-30,-21,17,-1,5,-26,-28,-14,11,-73,-6,0,12,23,-28,12,15,-19,25,8,0,-19,8,-42,35,-16,16,-5,-10,-10,42,-7,-41,12,15,-18,5,9,24,-14,-46,-14,41,-20,-3,-9,1,47,13,-3,8,-9,0,-28,1,17,-4,-25,1,19,21,-13,0,5,-18,15,-49,5,-1,-36,-33,4,16,-8,-38,2,2,-8,-37,-6,7,-37,-9,27,39,-8,8,6,-33,24,-31,-9,14,0,-47,16,1,-27,-10,20,6,-48,5,-4),
	(-57,-5,0,-22,65,-19,14,50,1,-4,5,19,15,-18,21,2,-15,21,19,-11,-31,-35,8,2,-39,17,16,-7,1,-51,-42,-7,1,-39,11,-10,-4,-3,1,13,28,-30,9,-6,11,-21,2,-45,4,-15,-1,7,5,2,2,13,-42,15,16,-7,-4,30,25,-34,-60,8,8,-10,-30,-19,-1,20,3,-14,0,-16,-14,-16,-4,-9,-10,-5,6,15,-24,-14,-10,2,-3,-8,-40,10,26,-14,-9,-25,26,25,-67,-19,-29,-13,-22,5,-7,-28,-13,-5,19,-6,-7,16,5,0,-34,-16,25,8,-22,34,7,-40,7,16,-12,0,20,2),
	(-52,5,0,-12,62,-43,9,10,-7,-24,-3,21,-6,-17,17,14,-29,16,12,-3,-23,-41,-34,-16,-43,-7,4,-12,-7,-26,-12,-21,-2,-29,3,2,10,-16,3,-3,0,-15,5,7,1,5,5,-9,5,0,29,9,14,-2,12,-11,-9,-6,0,-16,-4,22,10,-8,-45,26,-16,-8,22,-20,-23,12,5,0,7,-7,10,2,33,3,-15,10,-29,38,-8,-4,27,9,-14,-8,-30,7,44,-17,24,-59,35,46,-41,15,-27,8,-19,-31,-24,-10,-7,20,41,-4,10,-2,11,0,-24,-38,7,-6,-40,14,21,-9,-4,15,16,2,16,-1),
	(-67,14,-17,-1,8,-21,-3,36,-6,-10,-15,-3,13,-15,31,-2,-1,-8,1,14,-32,-32,-10,-38,-33,8,46,14,-13,-2,-11,24,-1,-4,24,14,13,-12,0,-6,8,-12,-7,-19,13,0,-12,-14,37,19,1,17,-28,-2,29,12,8,3,1,13,6,7,8,-25,-51,-8,-10,-5,3,-54,-4,28,0,-7,18,8,-9,30,12,22,-47,17,-26,40,4,12,27,4,4,-2,-28,-6,26,-32,14,-21,43,70,-16,-10,-42,3,-34,0,-14,-21,19,-8,28,-21,-15,11,18,26,0,-42,1,-11,-30,37,7,-19,32,3,2,-3,1,0),
	(-47,27,-3,-24,-42,-51,10,12,22,-4,1,25,14,-21,-10,35,-11,16,-2,-1,-17,-42,-24,-28,-24,13,31,22,2,13,2,13,0,10,16,20,-7,-14,4,0,8,-14,3,-24,12,0,-23,-1,27,11,19,-12,20,29,15,2,-1,19,-2,-15,-23,34,29,-17,-72,12,-34,-23,-6,6,-1,34,14,19,28,0,-8,13,-4,18,-20,18,-24,35,19,-18,17,24,-14,10,7,8,11,-37,-1,-12,31,12,-42,-5,-12,-14,-34,-4,-11,6,16,-4,27,-10,3,36,-11,5,9,-23,1,5,23,15,27,-5,13,-5,-15,0,23,1),
	(-40,14,-34,-16,-100,-11,14,16,13,-11,-16,6,3,-4,13,1,-16,9,13,25,-1,-12,-18,12,-6,17,-12,22,3,5,28,-7,23,-1,-16,-3,13,-26,39,-17,-14,-6,19,6,-12,12,-24,25,2,-15,1,-17,23,45,27,-22,11,18,25,-19,-2,28,26,-23,-47,29,-20,-22,-6,-1,16,0,-2,1,8,-1,18,11,-2,6,-8,15,-8,9,1,1,5,10,-26,37,36,31,34,-32,28,-1,20,14,16,3,-22,29,-32,-3,9,-22,14,17,17,0,-5,11,3,20,10,-57,-9,16,13,35,-4,16,21,2,0,8,-9,-4),
	(-41,7,-23,-6,-123,-14,14,11,25,8,-8,22,29,-26,22,20,-34,17,16,-8,-28,-29,2,-9,-12,8,-13,37,9,11,5,3,15,5,-3,22,1,9,25,-5,14,10,16,-10,0,19,-26,-3,6,13,36,9,32,16,-8,-14,22,33,6,0,-43,30,38,-29,-19,21,-30,-14,4,13,15,-11,-32,-5,20,-20,11,27,8,14,-26,2,-25,-19,4,-1,-4,-27,3,-6,17,22,14,-14,16,9,16,5,4,12,-34,-11,-37,0,-7,-13,11,6,6,-6,7,37,12,20,15,-48,-12,-1,23,21,37,7,32,-5,-33,24,22,21),
	(-38,-9,-14,0,-108,-15,13,12,8,0,-9,2,16,-29,4,9,-19,20,-30,10,-18,-18,-15,12,7,11,-55,32,-9,44,-7,6,30,7,-2,18,-4,6,28,-22,0,2,22,-1,15,4,-4,-33,9,-17,-1,4,24,36,4,0,2,14,21,5,-25,38,15,-30,12,-4,-6,-18,1,-7,-14,11,-47,6,8,24,-12,50,-10,-10,4,9,-26,-54,17,-8,-22,4,-20,18,15,22,33,3,11,16,25,10,44,7,-18,0,-23,0,16,10,-4,-9,-24,13,14,7,-19,-8,0,-50,12,5,-4,38,3,18,7,-26,-24,45,14,18),
	(8,16,11,23,-54,-4,22,-6,-4,5,-5,-4,43,3,-25,7,-38,35,-26,28,-37,-29,-27,24,-3,13,-72,30,-11,8,-5,14,22,37,-24,9,20,26,0,4,2,-1,-2,22,21,7,-18,-34,8,-2,3,-7,4,33,2,19,8,14,-5,-13,-28,44,40,-37,24,14,27,-17,5,2,-20,4,-30,30,22,-11,0,58,7,0,5,2,-29,-53,12,1,-2,-16,5,8,22,29,15,27,6,42,-14,-9,35,0,2,-17,16,-11,-11,-9,-3,-6,-1,-3,8,20,14,0,0,-33,7,22,10,9,-7,4,-2,-54,-34,56,6,15),
	(0,-2,-10,22,8,-4,4,23,21,-5,9,1,42,-31,-2,-4,-43,14,19,-7,-68,-36,-17,-4,-1,7,-44,51,-27,4,8,2,30,29,-6,-10,-2,-1,-41,-3,7,29,0,16,7,10,17,-22,3,-16,-9,-4,13,23,0,-12,8,3,17,-14,5,22,36,7,-6,6,9,10,27,-51,9,9,-52,6,5,10,25,50,-13,-23,0,-3,-26,-29,-7,3,-1,5,-10,17,2,6,2,18,17,31,-17,12,11,-4,3,-42,22,19,4,-2,20,13,-44,6,-17,22,24,-5,-11,9,-8,-6,-1,25,3,-22,10,-25,-16,41,23,17),
	(-3,-15,-4,25,59,-24,6,-26,2,0,-25,2,37,-5,15,18,-40,13,0,0,-65,-12,0,-9,10,21,-53,64,-10,-5,12,1,9,25,-10,8,-11,-15,-16,-10,1,23,-5,6,0,-8,-23,-23,13,-9,3,-9,-7,0,24,6,-13,7,4,-13,7,15,28,5,6,19,-17,10,8,-65,10,-12,-18,40,14,8,18,57,-13,-2,-24,27,-16,-3,9,-4,-9,-11,1,2,-25,26,-15,18,20,34,10,-8,9,8,-6,-26,33,-13,-21,-20,7,32,-22,-9,-14,12,8,0,4,53,13,-18,-10,1,0,-7,-12,-13,1,49,8,10),
	(22,-37,2,48,65,2,32,-49,-4,-26,-14,-12,36,-9,-10,12,-25,1,9,7,-37,-13,-1,2,-10,-1,-51,14,-11,7,3,6,38,36,-25,-18,9,-15,-25,-10,-10,7,-49,14,10,-20,-7,-47,7,25,0,8,2,3,-7,5,15,24,34,-1,20,31,15,-11,25,8,-2,-24,5,-40,20,-7,-37,17,-2,9,9,44,20,-24,-12,-5,-27,8,12,-17,-12,8,-20,-10,-31,15,-50,-12,5,62,-24,15,-3,-9,-13,3,17,-9,-10,-6,19,28,7,0,18,-13,-3,-6,13,65,12,20,-28,1,7,18,20,15,-27,21,26,14),
	(41,-3,-21,31,38,-16,0,-23,-3,4,-17,-2,-1,-3,-3,0,-6,31,-8,14,-10,1,33,-3,8,0,-2,13,22,-2,29,-25,5,40,-5,-12,10,-20,-24,0,-3,-23,-79,-34,12,-6,-18,-37,19,5,10,-5,-13,5,24,1,12,16,8,-16,42,7,8,1,4,0,-5,-26,0,-25,-9,24,-18,-5,8,15,-2,54,-25,-31,1,5,10,4,11,-13,-6,21,-5,-12,-35,20,-83,9,1,28,-8,0,-4,-12,0,5,25,-5,-5,4,8,0,2,-10,10,-12,-24,-21,6,69,-11,0,-39,1,42,-8,6,13,-23,21,17,19),
	(43,12,11,29,6,-14,-2,9,1,-26,7,12,12,-11,-7,-14,21,4,12,-8,-13,-6,19,24,1,19,12,-11,22,-3,20,-15,27,20,8,-10,17,-26,-28,22,-9,-15,-60,-19,21,-18,-41,-32,0,7,-27,16,8,-18,2,40,18,-16,20,-7,48,23,6,14,-33,33,0,-2,13,-8,20,19,-3,-52,18,2,13,-5,-11,-19,3,12,5,18,-3,-31,0,26,-12,-48,-32,37,-98,-44,-29,43,-35,-4,-25,22,-24,17,33,28,-5,6,-1,-17,6,-28,16,14,-16,9,0,12,-7,19,-6,10,27,9,16,-7,-35,-8,4,7),
	(60,10,7,-11,23,-2,-7,29,-29,-25,13,-19,3,11,-3,-17,10,26,1,0,-19,-8,55,27,-4,0,-5,-18,15,-4,0,-39,-18,39,-21,15,-7,2,-13,9,7,5,-51,-8,-8,-11,-5,-28,0,3,-25,-12,3,-16,-17,0,18,1,6,-2,30,-12,-16,18,-35,-6,20,6,1,-28,-14,-11,7,-51,-2,-19,24,11,6,3,20,-15,2,9,27,-33,-5,22,-9,-37,-39,2,-105,-32,-13,20,-64,-15,-8,39,-16,-19,42,32,15,9,10,3,-8,2,-11,14,-10,0,17,-4,-4,-1,9,-1,28,-14,-18,19,-35,5,32,1),
	(27,-2,18,-2,-9,-11,-13,11,-13,-8,20,11,15,8,-9,-2,9,-7,20,-6,10,33,32,28,8,-23,-8,-18,4,6,-21,-21,-19,32,-9,12,0,0,-11,-2,0,9,-23,-18,-22,-1,-4,-36,-18,8,9,-6,3,-28,-12,-7,2,8,33,7,17,-2,0,0,-31,19,-16,-8,6,-13,9,10,-6,-51,-22,-14,-19,22,4,3,-13,0,23,7,24,13,20,16,15,-63,-4,16,-101,-7,10,-3,-59,-46,-24,45,-10,-14,0,-1,8,6,1,-20,0,-17,10,11,4,-10,-16,37,5,4,-1,16,32,-11,6,25,6,-29,15,-2),
	(22,-15,-2,2,-28,-10,-9,16,-33,0,0,2,16,24,-45,12,37,6,-14,14,-1,46,14,7,25,-8,3,-48,-45,2,-16,-42,-3,31,-6,-20,14,-12,-1,19,14,-3,-2,-23,-10,8,-37,-30,17,2,36,12,-6,-30,-13,19,-16,19,-5,9,17,23,-5,-11,-52,12,11,7,-1,8,-9,18,-6,-54,-2,-28,14,-8,4,9,30,-25,1,15,-12,-4,13,4,-17,-45,4,-1,-96,-15,-8,-33,-61,-43,-32,10,-27,30,0,10,4,-9,-9,-14,-12,0,-19,-3,17,0,-8,2,-18,23,-1,0,51,25,-49,-41,3,0,21,6),
	(9,4,-15,-32,-7,28,-44,33,-52,-14,27,11,-1,14,-27,1,28,-7,-6,-7,-27,4,3,2,14,-25,30,-19,-43,-9,-4,-27,-31,-2,2,1,-6,-13,3,6,-22,16,5,-7,14,-4,2,8,28,11,14,39,-28,-8,-18,18,23,-27,0,1,-6,-5,-56,24,-60,17,-10,15,15,2,8,-3,-5,-40,1,1,-9,-10,11,31,16,0,-7,0,-9,3,-3,-2,3,-1,26,26,-88,-39,-7,-11,-35,-42,-13,14,-5,33,-4,36,-15,9,-13,-7,-9,-2,-14,-23,10,15,43,-4,-16,-9,10,-1,40,-16,-41,-7,-1,-4,-8,3),
	(37,-25,14,-56,9,4,-30,-15,-46,-10,-12,49,2,-19,-14,-13,1,-15,7,-38,-31,-4,-39,-1,7,-14,8,-46,-24,35,4,-19,-23,43,17,-14,5,15,4,12,22,55,4,-35,37,-14,0,6,21,6,-39,22,-24,3,-2,-17,36,-29,-10,-7,-5,-18,-107,-15,-7,-4,15,37,34,-8,-5,-6,21,-32,14,-16,0,-34,-20,-10,6,23,-18,-24,-11,-17,13,32,-17,1,36,0,-41,-52,-8,-29,-22,9,29,22,-4,19,16,14,0,-1,-16,-11,-3,-38,-1,-5,61,19,15,-18,0,33,-11,-8,36,11,-48,-5,-22,-3,29,24),
	(68,-30,18,-25,7,1,-31,0,3,-50,-34,60,15,-38,-39,-17,-8,4,20,-22,-17,-36,-29,-7,31,5,10,-7,12,16,47,-9,-9,37,49,6,19,29,-18,11,47,47,10,-25,44,-9,7,33,24,34,-39,10,-28,40,-1,-20,51,-53,-42,-6,20,-20,-82,-15,-59,6,25,16,5,-8,13,16,4,-18,0,-5,37,-27,-22,0,-12,36,-23,-42,-14,-24,61,35,-26,-7,17,1,-22,-58,-29,8,0,27,24,7,53,29,-15,8,-9,-15,-15,-35,-16,-35,18,-10,32,-3,0,-22,1,42,-22,38,87,6,12,-48,-21,-4,54,-16),
	(23,11,31,-5,18,-1,-11,-8,-8,-29,-18,15,-14,-1,-13,4,-6,4,9,-13,0,-3,-46,-31,1,0,19,-26,1,23,4,0,9,33,8,0,23,5,8,33,11,26,-3,11,30,-1,-9,-7,37,9,-51,-8,-15,12,-14,1,26,-13,-39,15,13,-4,-18,-2,-25,10,6,19,-6,28,5,-7,3,0,-9,-6,34,-37,-15,2,32,30,-14,13,-1,-15,23,45,-16,-5,-6,-15,0,-52,-6,-11,-2,-12,9,21,41,17,3,-26,-3,3,0,-5,-11,-30,-8,-5,10,5,3,-9,10,14,20,34,34,2,-10,-33,2,2,8,25),
	(3,-5,21,-15,0,2,17,-18,-26,-40,-6,20,3,-30,2,-3,0,-21,-22,-19,-13,-3,-23,-43,-16,41,-30,10,18,5,8,-22,-28,24,8,0,-5,-14,-29,9,-13,12,-2,8,-5,-3,13,7,6,2,-16,-32,3,38,-22,6,-1,-10,-27,-12,-24,-35,-5,15,-9,-29,-19,37,3,-18,10,-15,13,-16,-17,-16,13,15,25,11,-4,11,20,26,-21,-49,0,-13,9,-2,-21,4,20,-6,1,-12,12,2,-6,10,30,18,23,-24,-3,-3,-22,-1,-9,-9,-24,-11,28,1,-3,21,18,31,-16,45,7,-3,16,15,-1,7,-3,-20),
	(13,-11,4,-4,-11,0,18,-13,17,-10,13,-20,-3,20,13,14,7,-12,5,-9,4,-15,8,-18,14,-10,16,-19,-13,6,-16,-19,-7,18,-13,-10,11,15,-14,-19,11,-17,0,-7,-17,-19,-4,-1,1,-18,0,0,-1,-2,-15,13,-13,-17,4,18,4,-6,13,8,-7,15,8,-3,-2,-1,4,-19,9,-1,-16,-14,16,1,8,-11,10,13,18,-7,-2,-19,-7,16,14,1,1,12,7,-16,-3,10,-7,-3,10,9,17,15,0,19,-14,13,-10,-4,4,20,2,-18,-3,12,-8,8,-1,-8,-8,-20,-11,-10,15,-16,18,-11,-16,9),
	(-37,-11,-21,10,15,-6,-15,-21,30,45,17,17,20,-19,-2,18,29,19,13,19,-21,14,11,-31,-6,-6,0,9,23,8,-26,32,28,-45,-4,-11,-13,-1,-9,32,7,-26,23,-18,-25,34,21,-17,28,28,24,-4,3,-7,25,8,-9,15,5,8,37,35,37,-24,-30,-4,-44,11,23,8,21,32,-4,36,13,6,-28,35,-9,13,-38,-9,-26,34,26,-7,12,0,-12,-4,-20,-2,5,0,1,-24,16,13,14,51,-3,5,7,-9,5,3,-10,5,1,-28,-11,-35,6,35,22,-5,25,36,-38,1,14,-2,-7,10,6,-27,-6,4),
	(4,-32,12,-7,-37,-35,-4,-16,20,0,-31,4,22,13,27,16,-8,1,21,45,9,27,-25,10,25,-17,-35,4,2,7,9,-7,-16,-21,12,-15,48,-6,-19,10,-11,-27,40,-38,-27,-12,9,-18,15,6,7,-26,-3,4,55,33,-25,11,17,-9,1,37,-9,-4,-32,51,-9,-4,22,17,-25,-7,-19,14,-3,7,-12,18,20,43,-48,-31,-21,29,-22,21,44,-19,-7,14,9,-13,58,-5,21,0,24,1,-9,27,-1,-22,-17,-30,-12,-35,12,40,9,31,-4,-9,-28,19,40,-9,-7,19,20,3,25,9,-18,50,1,-22,33,-13),
	(-12,-29,26,-17,23,-10,9,7,31,12,17,-45,8,16,33,-1,36,-9,34,29,17,15,28,-13,20,-27,1,8,63,-6,-28,1,16,-36,-7,4,-2,-4,-16,32,7,-45,17,5,-9,28,14,-28,2,-22,11,1,-25,14,41,19,-21,15,26,14,-7,5,4,0,-7,0,1,-6,4,2,4,11,29,57,-26,10,0,0,12,40,-31,-27,12,47,3,13,34,-1,-21,1,-32,-28,-12,-9,16,16,-8,19,-15,20,1,-38,-26,-28,14,-23,5,1,-26,9,17,-23,-3,4,11,-3,3,6,-24,30,16,-19,-28,53,-11,-47,6,0),
	(-32,-17,-10,8,27,8,-17,9,47,39,7,2,24,-11,17,19,56,1,28,9,-1,52,0,-2,4,4,-12,-2,41,7,-60,-1,-7,-55,-45,6,-32,2,-5,0,-28,-41,36,19,24,-1,56,-83,6,-15,44,25,-15,-29,3,1,-44,20,-38,17,-23,5,4,-18,-1,-26,30,18,38,10,2,4,35,35,31,8,-30,14,-5,45,-24,-37,34,-13,4,23,0,34,7,9,-8,-27,-12,6,-26,-23,13,19,-6,-28,-19,-32,-26,14,20,14,-10,20,15,-4,-5,15,43,41,-33,16,6,15,-50,19,-15,-5,-30,39,0,-52,0,-11),
	(-42,-6,-9,-19,68,-15,-32,29,21,18,-3,14,-29,-31,8,7,39,18,33,17,-23,4,18,-17,-20,-20,55,-19,46,-31,-43,-10,23,-20,-12,15,14,36,-7,21,-12,-44,10,-7,0,2,32,-40,36,-10,17,45,-20,-50,10,-17,-47,-7,-23,-3,-6,-4,21,0,-25,-13,9,-12,7,-17,-28,2,5,-8,0,32,-3,-6,-7,10,-16,-23,-3,-57,17,12,46,53,-28,-10,-1,-20,-2,-4,-12,-48,7,9,-36,-17,-25,-26,-38,-8,-19,15,-22,-11,-22,24,-23,-1,10,6,12,-23,22,12,-40,5,-24,-38,-10,14,31,-47,14,-12),
	(-80,0,-5,-27,29,-17,0,29,19,-2,-12,17,11,-24,10,4,17,20,48,14,8,-6,4,22,-3,-18,26,10,41,-20,-39,-17,9,-37,5,22,33,12,-9,0,16,-43,8,0,-9,-4,9,-41,43,19,29,28,-1,15,20,-5,-23,9,27,0,-9,13,20,-39,-49,6,-26,-30,4,13,-32,-9,0,9,-14,16,-25,-10,12,0,-21,-32,-26,-47,-3,29,37,-7,-43,30,-40,-9,-17,-16,-12,-17,13,16,-22,-27,-28,-20,-41,-17,-26,-15,10,36,-5,7,24,5,-30,3,-9,-30,-3,-1,-40,28,12,-32,3,5,4,-43,44,-5),
	(-36,7,-3,-9,35,-20,-14,19,25,1,0,51,7,-37,30,2,-8,31,4,19,-17,8,-19,6,-31,-13,12,-25,1,-34,-30,-10,-7,-32,-4,-4,15,14,-21,24,0,-38,12,18,-8,14,14,-25,27,-12,10,-14,15,17,6,-4,-45,16,8,-6,-5,23,20,-16,-58,15,2,-15,7,9,-29,-5,-14,7,11,-19,13,10,13,10,-34,-14,-48,6,10,-27,34,-11,-20,-4,-48,-21,33,-3,-5,-33,-7,23,-29,-24,-56,15,-24,-4,-6,-6,-17,18,22,-14,-5,-11,-2,22,17,-42,-3,8,-50,45,17,-17,-9,5,0,-42,9,4),
	(-40,-14,0,2,20,-32,0,49,4,-25,7,18,22,-4,16,25,-29,0,-17,13,-26,0,-36,-50,-4,8,17,24,-24,-27,-4,-14,4,-37,0,23,22,-9,4,17,18,-11,9,-10,14,-23,-30,2,26,6,-10,11,-12,47,8,-9,-7,21,-15,-13,-3,17,-7,-1,-19,-10,-27,-14,8,-26,-8,-1,-35,-27,13,10,24,18,11,9,-23,4,-29,-7,12,-19,12,10,-3,-23,-12,-10,33,-51,-1,-48,36,55,-25,-5,-25,33,-19,11,-20,-15,14,13,-11,-13,6,5,5,4,3,-36,23,-10,-28,49,19,-22,19,22,-23,-19,13,-2),
	(-58,-7,-2,-6,33,-33,-1,31,15,6,-27,25,24,12,13,20,-6,14,18,0,-36,-27,-12,-28,-2,-24,13,-1,-10,-6,-22,-7,14,0,5,-10,16,-24,0,-14,6,16,-1,-15,-13,-19,-9,24,22,29,27,6,2,38,21,7,7,-11,-2,2,-28,23,16,-17,-21,24,-42,-18,14,20,-18,24,-28,-2,-7,10,1,2,-5,22,-31,-3,-12,40,1,7,-5,1,-2,18,-3,-12,17,-7,32,-53,27,16,-22,-29,-33,29,-20,0,-28,-4,4,-3,5,10,-11,20,17,-4,2,-29,-4,2,-14,10,8,4,13,-3,5,17,40,19),
	(-55,19,13,-14,-35,-11,3,6,5,14,-21,43,38,-31,9,19,-2,15,-9,23,-6,4,-12,-1,13,11,29,18,11,-14,12,8,16,8,12,-3,13,-11,31,1,6,1,15,-22,17,-9,-14,5,6,-15,32,6,15,37,20,-6,29,-6,20,11,2,23,30,-20,-44,33,-58,-21,20,15,9,13,-28,16,-5,-12,-10,2,0,14,2,12,2,58,-10,-20,10,6,1,-13,31,-7,27,-13,-5,-9,12,10,-29,-28,-36,36,-56,-19,16,-15,1,20,13,-9,-5,0,11,-11,-6,-34,1,23,9,15,19,19,-15,-2,13,41,17,14),
	(-8,32,-14,-5,-82,-23,19,-8,-8,24,3,4,21,-7,-3,15,12,7,-10,17,-18,-4,2,-2,10,-15,2,13,0,5,-6,-20,13,-5,-15,-19,3,-17,33,-13,8,16,17,10,-6,-12,-26,4,0,19,15,1,-2,24,20,-5,13,-5,9,-6,-45,17,9,3,-11,-1,-53,7,22,30,-20,16,-24,-20,-8,6,16,19,0,20,-11,20,-18,36,-7,12,0,6,11,-1,18,5,-5,-11,-10,-5,7,14,-11,8,0,-3,-40,6,23,15,4,4,-5,-7,-3,28,2,-6,5,-26,8,19,34,25,34,16,13,-4,1,44,15,24),
	(-35,35,-5,12,-92,-8,6,10,-7,-6,-24,8,37,-12,14,34,-19,9,5,17,-3,-16,19,14,18,17,-9,36,0,9,2,5,-10,23,5,-6,25,-14,15,7,-4,14,9,-16,-8,-13,2,-9,-11,3,18,-28,13,47,12,-1,24,15,25,-13,-17,0,19,-27,0,-5,-24,0,21,23,9,33,-51,-5,17,10,2,13,-14,7,-1,20,-24,1,25,-14,-20,-35,-5,-6,12,1,-7,-21,28,-12,-30,9,-1,12,-29,-11,-13,-16,17,-12,0,-5,12,4,23,31,3,4,-1,-40,0,8,4,42,45,10,27,3,-11,30,8,13),
	(-3,34,17,14,-101,0,18,-1,13,0,23,-2,39,-1,23,11,0,4,-14,15,25,-12,8,-1,30,-1,-35,23,-12,2,10,14,18,27,5,16,1,-7,18,-6,-7,10,36,21,13,15,-30,-33,-4,-7,22,13,19,55,13,5,8,2,17,12,-9,38,32,-17,10,5,-11,0,37,19,18,4,-28,21,2,8,22,17,20,8,12,4,-24,-5,-6,12,-13,-26,14,-2,6,2,-38,16,28,1,-7,29,21,-19,-8,-11,-16,19,-1,-24,-5,-6,-26,9,13,14,4,-25,22,-23,18,-1,8,23,36,-15,25,-50,-35,29,44,10),
	(20,-18,2,-4,-29,12,2,-11,-21,26,7,1,56,14,1,45,-23,0,-23,28,-4,-47,-11,-1,-3,5,-55,54,-26,39,24,18,35,27,0,3,4,25,-11,-15,7,8,24,7,18,27,8,-21,0,-46,-23,-16,2,48,20,13,20,10,9,7,12,44,8,12,37,8,-4,15,25,-25,3,12,-21,11,17,7,16,35,1,-18,22,29,-20,-37,15,-4,-4,-19,1,17,16,14,-64,28,7,37,-23,18,37,13,-2,-33,8,10,-26,-6,19,14,-27,-11,-4,13,13,-2,-16,-22,23,19,11,43,46,-27,15,-18,-36,34,40,31),
	(30,-1,1,15,39,-12,31,3,-14,-22,-15,2,20,13,-11,0,-34,29,-2,-19,-4,-55,-38,18,29,14,-54,41,-44,8,-4,33,8,37,-19,-17,13,0,-39,-22,13,14,1,30,4,16,-12,-15,10,0,-17,-9,10,22,8,-11,4,12,15,1,21,27,41,17,4,28,25,-12,47,-25,11,13,-47,44,5,-11,-8,33,17,-19,15,24,-41,-26,13,8,-2,0,14,8,-3,1,-78,31,30,39,-6,23,15,18,-20,12,31,-8,-38,3,8,43,-40,-31,0,-9,-16,-16,13,24,19,4,8,10,17,-34,25,-31,-42,46,29,28),
	(31,-41,18,31,87,-17,30,-8,-4,-5,-9,13,-10,10,-9,29,-11,28,-1,-5,14,-42,-15,-6,11,11,-42,31,-26,22,12,-3,28,25,-30,1,5,-8,-20,-18,20,-1,-6,0,9,-1,-39,-40,-19,-4,-1,8,30,39,18,5,13,-3,16,-21,33,34,9,-17,31,33,24,-23,11,-58,-4,22,-19,24,-16,-2,23,49,9,-20,-21,22,-38,7,-13,-15,-6,9,-26,24,-46,-3,-82,37,21,49,-14,18,-8,0,-20,18,48,-5,-12,7,26,5,-4,10,3,11,-23,2,-9,23,-8,8,13,40,56,11,1,2,-17,36,38,5),
	(7,0,21,8,97,-28,5,-29,10,-9,-21,-2,-4,27,10,30,-8,23,3,-8,4,-33,40,13,9,7,-17,19,6,19,-12,0,-12,5,-9,-18,32,7,-4,-2,17,18,-37,11,-6,10,-14,-38,31,25,-20,-15,13,-15,22,13,9,19,14,12,38,30,20,-10,0,29,-2,-15,23,-42,-20,20,0,32,-18,-9,16,20,7,-16,12,-3,-4,35,3,20,-3,-6,-1,-11,-33,24,-87,17,12,34,-1,-14,-8,-43,8,-11,15,11,-3,-3,15,5,-2,-14,20,7,-13,5,-28,61,-23,9,2,30,38,18,-16,3,-9,-4,44,20),
	(16,11,8,11,46,-31,4,-6,-9,-14,-6,33,1,1,-16,0,1,39,27,21,12,-6,27,0,16,-24,-17,26,23,13,-1,-32,11,31,3,-13,0,-28,1,12,30,-11,-80,-7,-9,-22,-30,-34,23,17,8,-5,43,6,-1,-10,24,14,21,16,16,17,16,23,-1,35,26,-25,-4,-9,-15,22,15,1,-5,10,-13,34,6,3,-12,18,-16,24,17,-11,12,-6,-16,-24,-38,3,-90,0,26,3,-44,5,-30,-34,-13,17,45,-4,-2,-2,0,26,0,-4,33,-3,-12,-4,-11,52,4,0,-18,-8,46,23,-6,34,-15,-3,50,-8),
	(20,0,26,32,0,0,16,6,7,-15,0,32,-27,26,-24,20,41,11,24,0,21,-8,46,6,10,-20,-30,-12,55,20,-25,-24,-12,25,-2,4,2,-19,-15,0,4,-20,-88,-10,-6,-5,-10,0,27,29,-19,0,33,-22,-1,28,8,33,-1,1,36,11,37,9,-33,16,8,-8,5,16,10,31,0,-54,-4,-11,15,7,-17,0,3,7,0,55,12,-11,-10,-1,-3,-34,-37,12,-88,-16,14,0,-20,-23,-51,35,-22,-7,36,3,14,-2,4,9,21,-7,12,-3,-26,12,2,52,-10,-7,-10,-14,65,0,3,15,-36,-3,23,12),
	(31,1,10,18,10,8,3,29,-21,1,-3,7,9,30,12,10,27,28,24,22,-5,-3,63,10,5,-19,-4,-25,19,28,-9,-32,-11,25,5,13,33,3,-11,12,24,-9,-67,-34,-14,-22,-9,-4,8,-2,-4,1,-6,21,16,37,23,14,-6,-10,3,-1,1,5,-36,25,9,-18,-8,-4,13,23,0,-63,-9,16,9,20,10,-10,3,-24,4,50,-9,-19,30,-4,-15,-61,-4,20,-95,-28,-20,22,-74,-38,-28,48,-35,16,12,-22,10,-23,0,-9,21,-6,6,6,0,6,18,40,-3,5,11,-6,46,19,-10,21,-21,-2,32,2),
	(47,-17,8,18,-12,8,16,36,3,-30,23,9,-8,5,10,4,16,23,38,15,17,12,27,17,28,-3,-7,-5,-32,18,-9,-39,8,24,29,-15,31,5,13,4,9,-1,-22,4,-11,-39,-11,-20,7,-18,-11,-12,7,-3,10,19,-6,-11,0,-3,18,5,1,24,3,26,5,-26,0,5,0,23,6,-72,0,-12,2,24,13,-4,14,-8,17,29,7,1,9,11,1,-58,-4,15,-82,6,-21,-2,-46,-15,-42,22,-7,40,12,-23,-9,5,13,-1,-11,21,17,7,-16,-25,13,20,4,0,6,-21,40,17,21,1,-25,-28,50,9),
	(62,-17,-4,12,-6,-2,-4,33,-7,0,19,2,8,0,-19,12,9,17,39,3,19,45,23,9,23,9,4,-38,-68,35,-2,-23,-10,30,11,-28,9,-13,14,-9,-4,-5,-38,-6,-5,-2,-14,-13,3,-23,12,31,-6,-40,5,33,-2,-1,15,-20,16,33,-20,22,-39,-1,4,1,-19,-1,-23,18,23,-62,-14,-8,34,13,0,20,6,-7,10,3,5,-14,22,-15,-2,-41,-15,4,-62,-9,-15,-11,-45,-24,-18,41,3,33,17,18,4,19,9,-6,-10,17,-11,-17,13,0,31,1,-7,-20,4,-2,31,16,-15,9,-14,-16,29,-4),
	(41,-15,0,2,-13,4,-16,39,-20,-7,18,2,-9,-5,-27,21,0,13,14,-4,-7,45,11,22,27,-30,27,-47,-49,-3,-26,-23,-11,-6,3,-8,2,12,45,8,-12,-6,-22,-41,20,-34,5,-5,21,4,-9,21,7,-44,-23,0,17,3,3,-7,33,-9,-66,29,-44,12,43,-4,-29,-12,-2,19,30,-67,-48,-27,-10,-12,-19,15,43,-16,-5,26,21,-31,-27,14,12,-29,14,29,-39,-22,4,-29,-20,-61,-18,29,-7,10,11,22,2,29,9,-25,9,11,31,0,5,1,31,-13,-7,-37,22,-18,43,-8,-34,-8,-31,-43,30,-10),
	(23,44,24,-47,-35,-22,-5,-5,-41,9,-12,12,-46,-21,-20,-37,2,-23,16,-30,-34,-12,-23,8,20,-19,1,-56,-21,18,3,-41,17,3,3,-11,20,3,31,2,28,-1,-50,-58,29,-7,-2,8,26,0,5,34,-15,-29,-10,6,26,3,2,-14,19,-4,-69,-12,-26,18,-4,0,-3,7,-19,-25,10,-17,-26,8,11,-23,16,-4,17,3,16,-27,-33,-21,-11,9,16,-32,17,-1,-36,-12,1,-27,-43,-37,-10,43,25,24,-21,2,-3,14,0,-10,-8,-19,-4,-13,27,4,0,2,25,-11,-3,-30,4,10,-35,-15,0,-30,-5,-23),
	(50,10,22,-11,26,8,18,-39,-38,-20,-57,29,-30,-33,-26,-26,-63,-4,-15,-34,-33,19,-53,-17,20,1,11,-24,-16,17,41,-36,34,0,33,2,13,30,23,11,34,18,-15,-10,48,-29,-6,5,22,17,-30,26,-33,9,13,2,33,-38,-4,17,-3,-51,-50,1,10,20,-12,-11,-15,1,1,-7,-9,-13,-16,6,33,-39,-4,12,30,44,-1,-33,-13,-12,45,-8,-29,-28,24,-18,-5,-14,-14,-27,1,40,2,11,45,4,-23,13,-1,6,-21,-37,9,0,-16,10,27,-1,24,-27,17,44,2,30,11,42,2,-68,-13,-29,11,-16),
	(23,-3,47,-5,21,11,-23,-13,15,-16,-40,-4,-9,-8,0,3,-27,8,19,-17,-8,-32,-62,-33,-2,7,14,-8,-1,26,21,-10,-10,-3,17,12,7,38,18,3,34,27,15,0,67,6,15,-20,27,-11,-24,8,-22,24,-5,14,5,-33,-16,-19,-16,-30,-33,5,-24,3,-5,-14,-2,47,-23,-4,-3,-16,-1,-5,21,0,-11,-16,40,29,22,19,-13,3,38,48,-8,-24,36,-25,-4,-40,-14,14,3,-25,0,22,29,33,-34,-20,-1,-7,-20,-4,8,-16,-26,1,29,-8,20,-24,-3,26,10,48,13,37,-1,-39,-8,-3,-2,0),
	(49,-3,4,-7,37,28,21,1,-4,-24,-2,41,25,-30,-14,24,11,-5,-18,0,-13,8,-39,-1,-17,10,3,-4,3,-1,-10,11,-17,-6,25,-6,-20,-9,-15,-21,27,21,23,18,11,-27,30,4,24,27,-8,-22,-14,28,-20,-30,28,-28,0,9,8,-3,-5,-14,-25,-13,-24,24,-9,24,20,-19,0,-9,-11,21,-10,-22,-2,-9,-3,0,21,13,9,-62,24,-9,1,-20,-4,14,29,-57,26,22,-25,0,11,34,30,4,14,1,0,9,3,-6,-33,-16,9,2,37,-15,-12,8,33,46,1,21,-12,-27,1,-24,-9,-6,30,8),
	(-23,-11,-30,1,29,-30,31,2,-19,28,34,15,-47,-30,-30,-6,15,40,-32,28,-26,18,11,27,43,-41,6,-11,-16,16,-41,-1,14,18,6,9,-8,-35,-13,-36,5,-7,-6,25,-2,-42,-13,-3,-2,-4,37,32,30,7,-36,-22,-28,14,9,14,7,-17,38,31,13,46,40,-2,-11,49,-21,-18,7,9,-10,15,-43,9,-22,27,27,-18,2,-23,14,40,-8,4,-13,3,-9,-18,22,39,-9,-12,19,-37,10,-25,22,17,29,-3,13,30,-12,-44,3,12,-24,-11,42,-20,-22,8,4,-14,8,-10,15,10,-6,-40,26,-4,18,-33),
	(-9,-7,20,12,-27,-1,11,-34,34,14,28,-18,13,-2,-3,30,20,8,14,2,29,1,-15,-51,2,-25,-21,6,14,9,-4,-4,16,-7,31,-49,25,25,-7,-1,15,26,27,-22,-8,25,33,1,1,-3,26,-3,28,-6,27,17,-17,31,-2,13,9,1,22,-39,-39,14,-25,-24,-21,32,-10,21,6,17,-20,-1,-4,-15,10,4,-30,-5,-4,10,0,26,16,-3,-20,29,-9,5,53,13,-1,11,19,6,-13,9,-19,8,-11,-8,7,-23,-16,23,-20,19,4,8,-19,7,58,15,0,22,-24,20,6,-7,22,54,10,-34,23,-42),
	(-1,2,27,-38,15,3,-5,0,-9,-16,-23,-4,4,-4,37,12,30,17,7,42,-23,34,20,-13,20,-28,22,-22,17,-10,-7,-44,-37,-41,-12,-16,28,-22,-6,5,-26,0,2,-35,20,0,10,-9,45,-14,-19,17,-8,-38,7,27,-2,0,31,10,-22,8,2,19,-48,29,9,0,31,33,-39,-3,-36,-13,-29,-13,0,9,24,29,-9,-23,23,17,-30,54,-1,21,12,21,-24,-2,-17,20,12,-1,21,-7,-25,6,7,0,-19,-21,28,-23,5,-4,-3,39,16,-10,-18,29,25,-14,12,-1,9,-4,21,3,-8,11,31,-18,26,4),
	(-12,-37,20,-30,30,-17,-6,9,37,25,-15,-27,-4,21,27,9,40,21,29,42,20,13,40,24,-23,-7,33,-11,37,-21,-41,-1,-12,-30,4,4,-21,2,-17,23,-22,-7,24,4,7,24,15,-38,38,-7,50,0,-3,-13,23,0,-33,11,18,15,5,-1,7,0,2,4,9,5,11,-20,10,28,0,22,-25,-25,-20,-28,21,27,-29,-40,13,45,-8,0,25,-8,-13,0,-27,-24,-10,18,-7,-14,-2,-12,14,10,-19,-14,1,19,17,7,26,17,16,3,-3,-15,1,39,38,6,5,8,-17,16,-2,-11,-17,15,-9,-36,6,15),
	(-40,11,11,11,39,-17,-6,6,49,24,20,-21,37,11,31,-3,38,-18,13,44,4,27,11,-30,-22,28,15,0,21,-16,-34,15,-14,-43,-20,36,-3,25,-18,0,-49,-24,23,-6,-9,33,44,-87,20,-9,26,0,-15,-40,1,27,-48,-11,6,1,-18,-12,4,4,13,-26,0,-6,14,-10,17,14,14,34,9,26,-6,13,30,17,-17,2,7,-7,4,16,4,0,-8,16,-4,-37,11,0,-10,-36,4,27,11,-33,-14,-25,8,14,23,24,-7,12,-2,-12,-13,1,29,15,24,-1,8,-9,-19,7,0,-26,-2,38,-1,-72,-4,-22),
	(-49,-8,8,-9,33,2,-19,36,29,-19,-12,29,11,-9,32,-1,30,21,31,1,3,12,0,-6,2,-12,24,-19,11,-30,-25,-17,19,-40,2,26,5,12,-27,27,-15,-59,35,4,19,15,-1,-34,23,8,27,-10,-4,-4,-8,29,-31,0,7,16,-21,-37,-6,-6,-47,-17,-34,-33,25,6,-11,3,7,-7,19,28,19,-22,-4,4,-25,-15,-2,-29,-12,36,28,5,-16,-10,-21,-38,16,-17,5,-14,-6,5,-26,-17,-35,-12,-15,1,19,6,15,0,9,14,22,3,10,1,30,-12,-21,20,-22,1,-16,-18,-30,5,15,-32,25,-12),
	(-28,-7,5,-16,24,-17,9,23,20,0,-21,9,-1,-3,31,-11,6,-1,29,4,18,40,8,-4,-30,-10,6,-17,33,-12,-27,-21,4,-31,19,-2,1,2,-28,-7,7,-46,28,-4,17,-18,-15,-16,5,-1,13,-11,-14,15,3,8,-29,-7,18,0,-13,-30,19,-19,-77,29,-9,-7,-9,4,6,-26,2,21,0,-8,21,-10,33,10,9,-16,-19,-63,-17,16,11,0,-22,-2,-15,-6,9,-33,14,-39,-17,16,-33,2,-21,21,-15,-7,-3,-10,15,6,14,16,20,-4,-4,-2,45,-36,3,1,-16,-17,-5,-18,-19,31,-5,-11,0,12),
	(-61,16,-8,-20,45,-48,-1,-4,3,-15,7,14,6,9,3,-15,-20,2,38,-4,10,3,13,-16,-22,6,3,-16,21,-48,-24,-7,-1,-9,41,11,-4,11,-16,8,-11,-10,-6,-3,0,-3,-5,11,22,27,20,-33,-9,9,12,-1,-9,-3,-2,-19,-3,-23,-18,-1,-74,-5,-27,-29,9,16,9,11,-6,4,-9,-1,-18,-6,11,6,-10,1,-25,8,9,-24,18,0,-11,-17,-5,-14,8,0,6,-55,-19,13,-12,11,-28,19,-31,-4,-13,21,1,31,-8,-5,10,7,-1,29,49,-13,-14,20,-14,12,25,-15,12,36,0,-11,16,11),
	(-59,21,1,-9,29,-24,-9,-6,19,0,13,24,29,-8,20,7,-36,21,2,16,5,0,15,-35,10,-1,-12,30,0,-49,6,14,24,-13,0,21,8,-16,20,12,21,-12,18,-11,8,-3,-6,11,21,17,-7,-28,-5,23,15,24,-11,12,20,-19,-23,-6,6,0,-27,35,-38,0,26,17,13,-11,-50,-12,-14,18,-1,17,5,3,-16,-9,-43,-9,-20,4,18,-12,15,-3,-8,-6,21,-7,23,0,11,23,-36,-22,-13,19,-5,-18,-39,14,10,25,26,7,30,9,1,16,0,-41,-6,-11,-11,21,16,-12,10,22,-7,40,23,-6),
	(-53,35,18,-5,47,-9,-3,-6,10,11,-22,20,4,17,27,2,-4,36,0,25,-12,23,10,-45,22,-30,11,6,-9,-39,9,0,20,5,21,0,0,-23,20,1,3,-2,25,12,-23,-46,4,22,1,20,3,3,27,7,19,-9,-5,17,14,8,-31,-16,0,-2,-12,17,-35,-3,67,1,7,14,-56,-1,-10,21,0,-15,0,1,4,6,4,44,-15,9,-14,-23,17,-17,15,-12,6,-5,3,-36,-43,7,-49,-25,-16,26,-12,5,-19,0,29,19,21,15,17,-7,-15,11,27,-28,-4,-14,-1,32,28,-11,0,10,-16,32,25,18),
	(-22,17,13,8,-20,3,29,1,-9,8,0,14,60,-20,14,45,-5,23,22,0,-4,1,-1,2,7,-11,13,38,-9,-45,-13,1,19,2,-7,-11,8,-15,4,-18,-8,12,22,-4,1,-12,-2,31,-4,13,47,-22,6,34,1,1,10,19,9,-21,-34,15,19,0,15,12,-48,8,44,33,8,20,-20,-4,-10,-7,3,-7,4,1,-15,-18,-11,22,21,0,-9,0,-25,-23,17,27,4,-16,15,0,-25,-4,-47,6,-22,23,-23,-18,5,17,-7,16,-2,-10,7,16,-6,10,34,-4,-13,17,0,14,43,15,-17,-14,-21,15,21,-2),
	(-8,38,-11,-27,-70,-19,-8,-33,15,-17,7,26,50,-17,18,5,-9,9,17,11,-15,24,2,31,23,-6,15,10,-17,-7,-7,8,14,6,2,-15,5,10,6,24,0,-3,7,-8,19,-30,-1,31,-1,-9,10,-19,6,31,22,8,10,0,15,1,1,-4,-23,-8,-15,33,-30,5,66,5,-1,20,-40,0,-21,-4,14,-34,8,14,-17,19,0,37,-14,-3,-2,1,-11,-32,40,-13,-30,0,-2,5,-67,27,-40,9,-3,13,-2,-1,16,20,-14,1,20,15,-11,22,7,2,34,-31,-18,23,2,30,13,24,5,-17,-37,42,44,-6),
	(-11,32,3,-13,-82,-3,-25,-7,-3,29,17,-2,45,-18,20,26,-15,31,0,-7,6,8,0,36,17,-1,-15,4,-2,-8,-10,3,11,-1,-6,0,10,11,7,-8,36,4,29,-11,-7,-35,2,-7,17,-13,1,10,19,20,-14,9,-8,11,-5,-22,25,-37,6,1,1,24,-16,-7,57,17,13,46,-35,20,3,-4,-18,-48,16,5,22,-16,6,-8,-4,11,-3,-22,-5,-43,6,11,-59,-28,-9,7,-39,-4,15,-1,-15,-21,0,-7,21,-16,-7,18,3,-16,2,-3,1,-4,23,-8,7,13,-1,21,36,11,7,-25,-38,37,33,8),
	(4,-3,-1,-11,-63,-1,-10,34,17,11,30,4,48,-16,-16,34,-18,28,-5,20,15,-20,-8,14,31,17,-45,11,-5,1,-8,8,4,-4,10,-15,-10,19,20,-8,9,4,26,0,4,-4,-2,-47,-5,-18,29,-25,2,44,19,-7,4,-11,11,10,1,-17,-28,17,22,6,15,27,28,3,31,44,-39,11,22,-1,19,-15,-18,-14,10,0,-7,-8,20,-14,-18,-26,7,13,32,14,-67,25,-14,8,-26,-11,5,28,22,-39,-18,-8,19,14,14,17,-4,3,23,-4,10,9,9,-28,-16,16,-6,27,9,3,6,-18,-16,15,10,-8),
	(22,-2,0,-22,-1,3,8,-1,27,4,20,-18,17,-5,-8,49,-53,29,0,31,55,-17,-12,19,15,5,-72,26,-62,18,-3,-2,-8,22,3,-26,3,18,2,-25,39,0,22,36,18,18,4,-31,-11,-9,34,-22,-2,30,36,16,28,2,29,2,29,-14,-7,2,31,0,35,-10,53,4,12,47,-3,49,-14,-6,-14,11,-6,1,4,9,-18,-41,-11,15,-18,6,8,33,-5,3,-78,22,6,-6,18,10,44,14,-14,-35,-4,12,-21,14,16,-5,-38,10,-8,30,0,1,-4,-24,-16,27,-9,40,43,-14,-1,-18,-30,-9,24,14),
	(14,-15,27,10,49,-5,-10,0,20,3,15,-9,26,4,-16,23,-36,10,11,27,46,-15,-3,4,21,-20,-44,9,-33,0,0,-5,16,10,-15,-1,8,5,-10,17,25,3,29,38,7,28,-23,-40,19,-14,27,13,2,13,10,10,20,13,10,1,8,31,25,0,-4,-2,9,-15,23,-19,13,39,2,34,-15,4,5,16,6,0,1,14,-31,-1,8,3,-7,-26,-13,48,-9,-4,-79,51,25,2,27,-10,2,-16,16,4,22,-21,-26,4,20,0,-35,-11,-3,19,-28,4,-11,-13,-10,30,8,29,46,-23,-14,2,5,6,32,15),
	(26,-11,22,-5,74,-13,4,-25,20,-23,-23,19,0,9,-17,0,14,28,0,26,49,-23,30,0,30,-15,-38,23,-4,18,0,-14,18,-4,-18,9,22,-11,-7,1,28,-46,10,20,-8,2,2,-6,0,14,12,-9,10,16,29,-3,14,13,12,-15,14,2,32,-28,9,5,37,-15,20,-25,-17,16,47,51,-12,-22,-20,15,15,-6,-19,13,-12,18,-3,-13,-6,-34,21,-3,-47,22,-68,23,21,12,36,5,-12,-57,5,4,45,11,-6,0,12,-13,6,9,2,0,-25,-10,6,16,20,-1,26,33,52,-4,-20,4,-30,-13,27,19),
	(15,-24,29,36,63,0,-17,-36,16,-28,0,40,7,39,10,22,7,26,17,14,51,-42,31,-7,29,2,3,23,50,7,-10,-24,20,-21,-4,0,26,-14,0,8,10,-48,-2,5,-8,2,-8,-26,-3,3,4,11,48,-16,17,-35,-11,39,-1,-8,-2,16,19,-6,3,1,43,-2,23,3,2,31,64,38,-30,-17,-3,18,-13,10,-13,5,-25,47,-2,2,1,8,-2,-12,-35,7,-35,6,22,-17,23,-33,-46,-61,8,8,31,6,0,-6,6,-12,12,11,-4,-4,-11,9,-18,27,5,4,12,8,17,-4,1,-6,-9,-33,30,1),
	(9,-8,32,43,29,-5,20,0,18,-29,8,21,-21,35,-8,8,8,18,39,35,21,-8,65,29,11,-20,21,37,30,-13,-17,-11,15,-23,-3,0,27,-3,13,8,32,-24,-48,-31,-14,0,-23,-15,35,33,10,18,15,-11,14,0,-10,33,10,10,24,-2,42,-13,-5,5,26,-10,9,30,8,3,49,33,-34,-28,-27,25,6,-7,16,0,2,25,2,-15,-30,-10,-20,-30,-18,-1,-41,-26,51,-11,-35,-7,-65,-25,6,11,17,14,4,-10,21,-5,27,-7,8,-4,6,31,8,33,-15,-12,6,26,26,-1,-16,-6,-16,-35,10,31),
	(44,-7,11,19,-36,-6,10,0,9,-18,-11,25,0,0,-5,23,18,28,13,15,24,-29,40,18,-2,-6,8,10,51,23,-3,5,0,-26,-6,-4,28,10,10,7,-18,-59,-58,2,-1,-14,-29,-22,21,24,-24,20,9,-14,17,-12,21,28,10,17,38,-1,50,-15,-48,10,9,-5,18,14,-3,25,55,-34,-19,-15,-12,9,12,4,19,-10,-5,17,11,-9,-19,0,-6,-28,-9,1,-48,4,29,-18,-49,-37,-53,29,-8,-4,9,7,20,18,26,12,24,-33,-6,13,1,-3,-22,48,-22,-20,4,19,56,7,2,20,-35,-27,30,12),
	(27,9,1,31,-44,-9,1,19,10,-23,17,7,-12,0,18,2,-3,24,40,28,42,20,17,-14,22,-11,-5,1,13,11,-11,-7,12,-36,7,22,18,13,28,22,21,-62,-73,-10,18,-17,0,-27,0,7,0,22,30,-17,3,18,19,18,-9,-20,24,13,31,-13,-59,2,14,11,-19,6,7,37,9,-69,-47,-3,-6,-11,9,15,21,-12,16,36,-15,-14,17,12,-23,-32,-15,8,1,-17,-31,-1,-76,-31,-23,48,-16,6,16,10,22,14,21,-16,-16,-25,-9,15,-11,10,14,35,0,-8,4,-2,49,17,2,-4,-11,-37,12,9),
	(71,-7,9,31,-49,7,-5,8,-35,-2,-10,22,-11,-13,17,-18,1,28,15,7,20,37,25,-9,2,-2,32,3,-54,31,5,11,18,-12,12,2,14,8,43,20,0,-26,-58,-24,11,-18,-21,-11,-8,9,1,-11,28,-19,8,6,3,4,22,13,26,-27,4,16,-42,-1,33,-2,-34,19,14,13,17,-62,-27,0,-1,8,15,23,32,-13,15,5,-11,-6,-20,1,15,-82,16,5,-7,-7,-30,-5,-63,-6,-1,47,3,0,6,10,0,-17,-1,-2,-17,-12,11,1,-18,-12,20,6,-17,0,-11,-16,27,18,-25,4,-32,-7,3,-8),
	(29,-22,-5,22,-56,0,-8,20,-9,-10,14,0,-15,10,-19,12,7,41,54,34,35,29,26,-4,2,10,37,-14,-59,11,-19,-21,13,-21,17,-9,22,0,42,11,0,-41,-45,-38,2,-40,-14,-18,30,5,-9,33,-15,-19,6,24,15,17,21,-18,39,17,-29,1,3,-24,25,-19,-8,32,7,41,42,-82,-21,-18,-4,0,-5,12,-15,-1,-23,-1,14,2,-2,-19,-13,-32,-4,25,-16,5,-19,-2,-41,0,3,43,-19,-13,21,-7,3,-7,-2,8,-12,-21,-5,-25,11,-8,47,40,9,0,-2,21,18,-11,-19,18,1,-48,22,14),
	(46,-8,-8,-11,-28,-5,1,-4,0,2,34,-3,-15,-12,-19,15,-21,29,15,0,30,33,8,17,8,1,8,-29,-57,5,-18,-29,23,-26,13,-26,34,11,12,32,2,-15,-61,-46,-3,-16,-15,-17,41,-18,43,42,34,-40,-29,5,20,-15,24,17,19,15,-42,5,-18,0,27,-19,-18,28,0,33,40,-58,-57,-34,25,-1,4,24,-16,8,6,-1,-2,-26,12,-5,-27,-21,26,-16,-11,-1,-6,-30,-37,-11,-11,17,0,4,-13,25,41,6,-34,-8,-21,-19,12,-18,-2,9,18,4,-23,8,-2,-27,24,12,-29,9,-14,-25,29,-18),
	(72,27,39,-21,-43,-19,-9,4,-38,4,-17,11,-31,-21,-27,2,-61,15,2,-35,28,16,-21,23,22,-30,35,-51,-41,6,29,-51,-7,-4,8,-48,38,24,40,17,7,-2,-27,-25,12,-8,-32,-6,42,-38,6,40,6,-7,-3,24,46,-17,-18,-2,32,-24,-96,-8,7,70,26,-34,-9,37,-28,-11,52,-41,-77,-5,17,-33,9,-27,17,22,-16,-52,-3,-32,15,4,-8,-15,26,33,21,-36,-25,-48,-27,-31,24,-1,-9,15,-13,26,25,-8,26,-14,5,-6,33,-22,0,-22,50,-41,-19,14,25,3,-11,37,-34,-18,-35,-26,6,21),
	(47,26,55,-6,-37,-9,2,4,11,-8,-31,16,-23,-24,-31,-45,-43,-15,-21,-14,-2,-42,-43,7,28,-20,36,-52,-37,33,44,-70,-11,1,27,24,6,50,27,39,29,10,-17,-17,80,-17,-5,36,31,-52,-12,44,-24,15,-1,32,33,-42,-35,11,-5,-35,-59,-4,5,55,16,4,-39,10,-30,-4,16,-23,-15,10,47,-24,-13,-4,22,73,9,-52,-9,-1,10,30,-8,-39,8,-19,-6,-46,-16,-19,11,-3,10,31,60,9,-37,7,19,4,0,2,18,-15,37,10,17,18,17,-63,-25,-10,44,0,9,43,-27,-38,-33,-21,19,49),
	(-8,-15,9,0,-10,21,8,-16,26,-36,-2,16,27,-40,0,14,-47,3,12,0,-2,-32,-60,11,1,34,42,-26,-12,9,-2,-12,-13,4,39,25,-12,33,25,1,12,26,-4,-1,58,14,12,-2,39,-16,-10,22,-15,-5,12,21,35,-9,7,-1,7,9,-17,22,-61,-5,6,-9,0,33,3,30,-10,-16,5,10,45,7,-4,8,9,29,-10,-37,24,-36,1,39,9,-29,2,-11,6,-47,30,10,1,-23,-23,19,25,28,-12,34,37,21,36,23,-8,-18,30,7,27,-6,31,-22,-24,-8,54,25,11,1,-36,-35,-30,10,6,6),
	(11,-2,1,4,-8,-27,16,-2,10,-5,33,30,6,-16,-8,-12,3,17,27,0,48,15,-3,6,39,0,10,-37,-4,-2,41,7,0,9,45,6,0,-1,-10,-21,24,46,-29,-26,10,6,18,36,31,-6,13,34,21,-1,13,13,15,-15,16,3,7,4,-14,-7,-8,19,20,32,2,11,0,36,16,5,-16,-8,8,-21,-18,4,-5,20,4,-17,7,-22,-1,9,-17,-9,-17,34,23,-49,6,-5,-12,1,-5,-6,-1,34,-3,38,40,18,6,18,-42,-16,27,8,22,-2,11,-12,4,25,30,6,8,4,-15,-14,-3,-6,32,13),
	(8,-12,5,8,6,-29,12,-23,-5,25,0,-12,-6,13,7,-3,-21,-11,26,20,28,-11,-12,7,9,9,-4,18,-7,9,0,-2,15,-9,26,-23,28,-24,-14,6,0,-2,-7,0,-26,5,-10,-9,8,22,0,10,13,10,18,9,-9,13,8,1,0,5,-9,-23,3,10,-4,-1,-2,8,-1,-1,7,25,-9,0,9,12,32,-6,7,-20,-11,14,-11,-8,-5,-15,5,16,-10,-19,7,-12,21,8,-28,0,-1,15,-14,-6,-12,-28,18,-15,-11,9,-25,5,25,-6,-23,14,8,6,-16,15,-8,16,19,-5,-14,24,21,-2,0,0),
	(0,1,23,11,22,2,-8,-34,29,30,-9,-1,5,27,19,1,8,19,13,27,10,10,8,-23,17,4,18,0,20,35,-30,-1,-24,3,18,-38,26,0,-4,2,-6,37,31,5,-16,14,13,12,21,15,-13,-18,30,7,0,12,-5,8,7,13,28,15,-12,-4,-43,22,-18,-21,-18,41,-20,23,-13,16,-30,9,-4,2,-7,5,-20,-14,-24,37,-10,38,14,0,-2,-6,17,5,32,-22,13,8,3,-20,10,12,-30,-24,-3,-3,-5,-23,-12,-1,-15,18,5,-22,-15,-5,5,-32,-23,19,-22,1,18,-18,38,42,23,-35,22,5),
	(11,9,4,-26,4,-8,-10,-6,-17,-1,6,-3,-24,1,19,-27,10,-28,22,16,-23,15,32,10,0,-17,29,-15,14,-18,-27,5,12,-20,-5,26,-9,13,6,10,-21,-1,13,-9,-6,-14,12,-4,15,34,-4,2,12,-13,2,3,3,20,-4,5,-4,-8,-14,-7,-54,-17,-8,-11,29,-18,-14,12,-37,-16,-6,-17,12,-11,14,44,-18,-17,-22,20,14,21,-10,-13,10,10,-27,-11,-10,-13,-14,-1,-2,-22,-4,-24,14,-7,24,-2,28,0,-3,6,41,-14,4,-18,-7,19,36,-24,-17,10,1,-15,4,12,-18,-15,-4,-37,-28,-8),
	(3,5,-17,5,9,-21,-16,-29,41,-1,25,-17,8,9,-12,-1,10,2,9,27,17,9,14,-6,4,12,16,15,35,-29,-42,3,2,0,24,7,-1,-12,-21,-9,-4,-12,28,29,-10,8,35,-31,23,1,42,5,13,-20,0,22,-36,26,-2,1,-5,-5,-35,6,-23,4,9,3,4,-33,16,2,-24,29,-11,-13,0,23,7,16,-25,0,0,25,19,17,-5,-6,-4,25,-53,-41,-11,30,12,-20,25,-20,22,0,-9,-19,-7,5,14,27,-14,-13,25,10,-11,6,15,19,17,10,25,24,-21,10,18,-2,22,-6,9,-47,1,5),
	(-29,26,19,-4,4,-7,-15,11,2,29,14,10,12,18,0,-7,0,-18,6,4,-5,42,34,-36,-14,2,25,3,17,0,-31,38,-31,-5,-29,-6,-17,23,15,-1,2,-44,29,17,0,21,35,-77,0,10,1,0,3,-5,-7,-14,-47,11,8,13,-29,-15,-32,-21,10,3,-27,-26,19,-11,10,20,8,41,17,0,0,-16,13,-3,-29,-25,-37,-12,0,17,29,19,-19,32,-17,-48,12,-15,-15,-17,9,0,16,-34,0,-20,-4,-20,24,-3,-12,37,27,-19,-23,9,-5,0,14,19,8,42,-50,-2,14,-23,-21,16,5,-46,-1,-10),
	(-49,20,17,-22,26,-17,11,54,23,-20,11,-6,22,-7,11,5,-17,-8,10,-8,-16,3,-7,-32,5,-14,12,-6,7,-22,-10,-15,0,-46,-27,19,17,30,-3,14,8,-43,24,-7,18,-15,15,-37,0,7,-7,-25,-3,24,19,23,-74,-14,-11,-19,7,-41,-17,-24,-69,-3,-20,-27,8,-26,-14,-19,26,4,-11,16,-4,-21,31,-8,-35,16,-44,-39,-13,10,-13,-20,-37,-5,-36,-29,20,-14,13,-8,-25,31,-49,6,-33,-32,-8,1,15,12,18,21,-23,5,6,13,13,-5,18,-9,-5,34,-25,1,18,-11,-3,37,7,-37,-7,-20),
	(-57,32,-4,-25,-6,-32,27,-5,12,-50,0,10,11,5,3,-35,-45,3,7,11,-1,6,-16,-26,-14,-7,3,-16,-12,-16,3,-7,15,-11,-12,10,20,27,-15,14,7,-9,-14,2,9,6,4,-19,19,11,-17,-17,0,44,-9,16,-39,24,29,-15,-19,-45,-15,-19,-62,13,-38,-4,29,-23,18,11,-14,9,21,8,2,-25,19,11,7,-1,-35,-38,-13,-35,-3,-2,-15,5,-33,-9,23,-4,29,-17,-29,-1,-19,24,-43,30,-45,2,-8,19,16,16,27,-25,13,22,-11,17,20,-43,-2,-2,-22,-6,3,-7,-4,1,-22,-3,-12,15),
	(-74,10,6,2,21,-2,-15,-12,-1,-2,34,44,21,18,8,-3,-33,9,-1,-10,8,20,-6,-10,-16,10,9,-1,-12,-47,-20,7,-12,-23,14,16,-1,12,-16,-4,25,-25,30,-23,0,-5,11,7,12,16,-2,-16,0,24,13,2,-32,3,22,-9,-17,-46,-19,2,-38,27,-33,20,49,1,-1,14,-39,14,14,18,-32,-10,8,-33,9,3,-17,7,12,0,16,-7,-13,9,-36,12,12,-11,20,-9,-33,-18,-2,0,-14,7,-35,-6,-31,-7,23,15,10,2,10,6,19,22,26,-4,-13,-3,-25,36,-6,-18,1,13,-7,19,16,-5),
	(-42,-1,8,-22,57,-6,3,24,10,-20,38,16,17,20,21,0,-41,-2,21,-3,-21,13,2,-41,-8,6,19,26,-33,-11,13,0,-18,-9,6,-1,-11,-10,17,11,19,-15,7,0,7,-17,1,-15,8,18,-25,-14,-10,34,3,-9,11,13,25,-10,-20,-35,-15,-18,-11,7,-34,-13,50,4,-11,23,-31,-15,-5,27,-5,2,7,-14,-10,-1,-42,-3,25,-16,21,-14,3,-46,-29,22,11,-2,4,-24,-29,8,-22,21,-33,36,-27,-9,-14,12,20,30,2,-2,22,0,14,9,13,-6,11,27,0,40,5,-9,7,0,-14,14,25,1),
	(-26,9,10,-20,36,-16,-4,23,8,-18,29,37,40,12,16,12,-39,16,-8,-33,-14,-3,18,-42,-9,-8,15,9,-10,-39,-7,-2,-14,16,26,-2,-3,-34,-1,5,12,-12,37,12,-19,-26,7,4,-7,-2,-13,3,10,38,-15,24,3,4,18,-2,4,-44,-6,17,-5,18,-28,4,78,-5,-1,-8,-22,3,-26,-14,8,-23,17,3,-6,1,-3,45,8,-18,8,-5,-5,-60,1,21,36,-6,-1,23,-69,18,-38,4,-21,39,-14,15,0,-7,19,18,12,5,2,34,-16,8,8,3,7,12,15,-2,-5,-3,-1,-7,-28,11,20,10),
	(18,44,14,5,-9,-26,-18,-30,0,-14,40,31,32,8,20,7,-14,16,3,-32,13,9,22,-14,28,2,17,-13,-20,-32,-4,-12,-15,-7,-3,-3,-6,-26,-22,-11,36,-19,36,3,0,-31,-20,-11,8,10,-11,-1,-10,17,13,20,-6,-8,20,2,3,-33,-33,0,19,21,-80,23,55,13,-10,10,0,7,-17,5,12,-15,3,-26,3,13,19,7,2,12,29,-22,-23,-34,-4,18,6,9,19,27,-30,5,-66,8,-14,5,6,-11,6,-5,6,13,19,13,-17,27,-23,3,-4,7,3,-2,-7,6,11,16,7,7,-19,15,9,14),
	(15,35,13,-24,-53,12,-27,-12,3,8,33,21,35,-4,18,-13,-21,11,3,-15,13,16,-13,14,13,9,32,-40,-37,-20,25,17,-19,42,17,-4,1,-11,-6,-8,33,19,15,17,29,-49,-23,-11,4,-24,-23,10,-15,21,-10,-9,3,-3,5,-11,15,-86,-31,-22,12,31,-45,-15,65,37,14,1,-15,-18,7,-32,1,-16,-3,-27,-14,-3,10,18,-20,18,24,-29,-3,-35,1,-9,-17,-11,-16,9,-19,-3,-11,9,10,10,0,-16,31,-26,5,-15,18,17,-9,24,15,-12,15,-12,-4,32,16,-19,26,34,-2,22,-25,15,29,7),
	(9,24,4,-14,-77,10,-29,-13,-8,-2,42,1,17,-1,-8,11,-16,-22,17,1,48,16,-14,47,8,4,5,-28,-17,-12,-4,19,5,15,5,-19,14,0,15,32,45,-12,24,5,-1,-36,-20,-10,21,-47,6,14,-28,25,12,-5,11,-1,16,11,35,-75,-42,-18,-21,12,-9,-13,64,27,-14,1,-8,5,21,6,-4,-19,7,-3,-6,-14,0,-37,4,-1,1,4,18,-25,2,-12,-28,-15,-11,10,-11,9,-1,-3,-6,-34,14,-14,32,-22,-15,8,12,4,18,10,20,-15,14,-17,2,11,19,15,24,26,-3,18,0,0,8,1),
	(15,0,7,-15,-57,-1,0,30,16,48,50,10,26,4,-28,4,-36,9,22,9,67,-3,-3,46,0,3,-47,-8,-17,-7,-10,-3,-25,31,1,-8,22,32,-7,11,30,-8,5,-1,23,22,-13,-50,20,-30,13,-11,-30,39,32,15,25,6,-3,15,3,-111,-43,-5,17,-14,40,3,35,28,6,12,13,16,16,-27,-9,-37,0,8,37,6,-2,-92,-4,26,-41,-30,-17,31,29,-16,-54,9,8,-14,24,-7,11,4,-2,-68,-11,-11,41,20,32,20,8,9,28,-16,-2,-11,11,12,-8,46,0,23,22,12,-4,29,0,-13,9,-7),
	(11,-8,0,-4,10,17,-6,15,8,40,34,-40,25,-1,-11,15,-57,-14,7,14,50,0,-45,21,18,5,-56,2,-38,17,3,14,7,3,6,-22,5,0,-32,17,40,0,44,39,-11,26,5,-72,15,0,2,11,-14,39,4,14,5,39,31,-7,-6,-87,-31,-8,27,6,36,8,47,22,1,34,20,46,-9,6,1,-38,-8,-3,5,-8,-6,-76,-16,13,-46,-21,16,42,35,-9,-37,48,-18,-5,13,-18,38,-12,-15,-64,0,4,19,-4,10,-10,-9,-13,30,18,-10,-6,-20,-11,5,36,-7,31,-5,-28,19,11,-2,-11,9,-10),
	(-9,-38,33,-29,60,24,3,12,32,-9,28,-22,28,40,-17,17,-41,2,23,-6,69,-14,-57,12,-5,8,-62,20,-2,4,-16,-25,-6,-19,27,3,5,7,3,4,-6,-20,18,38,-6,42,-12,-56,-13,21,17,-25,22,41,43,0,-6,19,13,-16,2,-28,-14,0,32,-10,39,-20,10,3,0,21,29,54,-21,-6,-13,4,2,-9,-18,-28,-36,-9,-14,19,-40,-11,20,54,-33,-4,-28,56,30,-32,21,20,20,-39,15,-26,5,8,15,-6,37,-23,-2,-21,7,10,-21,-3,-13,1,-19,33,31,2,-4,-16,-4,9,9,-57,14,21),
	(1,-32,32,16,62,-21,-20,2,5,-11,5,15,-3,24,-26,29,19,-1,15,25,32,-30,1,-26,2,7,1,7,34,8,-20,-19,-3,-44,12,16,8,19,-12,6,-25,-50,7,21,3,18,-20,-10,16,19,22,-18,2,0,32,-5,-18,35,33,-7,4,21,38,-16,4,17,34,0,-8,5,20,7,67,51,-40,-3,-17,13,-1,17,-1,-6,-13,37,5,18,-21,2,0,2,-46,7,12,2,27,-38,47,-2,-36,-93,15,12,0,-10,6,11,6,-20,26,11,27,22,-12,18,-29,-6,5,29,12,15,-12,-7,0,5,22,-33,3,6),
	(-16,-4,21,7,53,0,-17,18,4,0,-19,7,9,27,0,8,7,-13,14,6,51,-22,58,4,6,7,17,8,47,-3,13,3,13,-72,24,5,-1,27,20,9,-13,-64,36,13,0,-25,9,-27,9,28,13,12,3,2,26,9,-5,13,20,13,35,22,53,11,-37,-1,22,-23,0,24,4,25,55,42,-37,-7,-15,21,7,24,-15,4,13,52,15,-3,-22,-6,-22,2,-41,15,43,-19,27,-33,38,-12,-28,-39,-11,-17,12,-14,23,-9,39,-13,26,0,6,6,-24,19,-12,-25,4,15,3,0,-6,13,-30,22,-23,-44,-11,29),
	(1,-10,20,33,-4,-1,-15,-8,23,-14,6,7,8,10,6,21,40,11,6,30,43,-25,50,-10,7,10,15,10,47,21,2,-25,27,-74,-18,22,31,6,16,31,4,-65,-11,12,11,-3,-5,-32,11,31,-5,-7,32,-8,29,4,-20,25,11,-15,2,6,47,18,-15,-6,40,-17,15,45,-11,-11,57,28,-56,-46,-11,0,7,0,23,-7,8,17,17,4,-22,-21,-33,-39,-28,-18,44,-46,40,-32,-21,-10,-54,16,14,-9,2,0,27,-4,31,1,43,-14,28,19,-4,10,-13,21,-15,1,14,13,-7,16,-31,26,-14,-56,12,6),
	(-6,-6,16,24,-40,-16,23,-4,-7,20,0,-11,8,23,-15,7,32,13,11,29,-2,-3,68,-15,16,0,15,29,28,18,5,10,14,-94,-11,21,8,7,19,3,-16,-69,-55,10,0,-13,-12,-15,6,49,5,11,27,-11,-19,6,3,24,26,-1,29,-25,42,9,-22,2,45,-17,-12,18,23,8,33,-12,-29,-21,0,27,-9,7,7,-11,-7,-2,-8,-24,-41,-4,-35,-40,-28,-17,47,-16,21,-26,-41,-17,-33,60,0,-18,19,-1,19,9,25,13,7,8,32,4,-12,2,7,14,-4,18,-5,-17,0,-13,-25,5,-19,-45,11,6),
	(-4,22,24,-3,-34,-9,28,-23,-10,2,-10,-15,-16,-4,8,-8,15,21,26,18,1,38,19,22,0,4,34,21,-9,2,-27,6,18,-87,-19,23,12,-11,20,22,-13,-58,-79,-44,-12,-39,-18,-23,8,40,23,3,23,-51,14,5,-33,39,35,-15,0,-23,10,0,-57,17,28,-20,-1,45,8,23,43,-46,-27,0,-7,-5,28,32,13,4,8,-10,3,-17,-35,-21,-35,-65,11,1,33,6,-22,2,-87,0,-12,72,-2,-22,31,18,19,4,26,28,-2,-8,30,-17,-15,0,10,50,8,19,-3,-23,-22,3,-41,7,7,-27,19,7),
	(44,-14,28,11,-55,0,-1,-18,11,12,9,-12,-23,-19,-3,-22,0,5,7,6,7,33,21,9,-26,3,20,-6,-58,14,5,5,0,-50,17,0,-3,-4,38,26,-18,-31,-60,-48,8,-27,-14,9,33,23,18,1,20,-27,-30,17,-2,2,23,-22,26,-4,-12,15,-40,9,21,-1,-51,40,8,3,45,-79,-34,-4,-5,-20,7,41,18,0,-3,-6,13,-24,-3,-15,-25,-66,12,4,32,-5,-26,-22,-66,-17,-20,88,10,-11,1,-11,30,19,10,39,5,-34,17,5,19,1,39,31,-8,-1,0,3,-17,-8,-6,16,0,-32,-1,4),
	(11,-13,28,19,-42,-26,-3,6,-21,21,1,-34,7,13,-13,2,-41,16,37,19,20,36,7,-14,-8,-11,10,-7,-45,38,0,0,2,-31,14,-15,3,-8,46,25,5,-39,-46,-36,26,-43,-3,-25,31,-3,27,14,19,-20,-3,22,-3,17,16,-6,32,-2,-14,3,3,-19,3,-33,-2,3,22,61,46,-91,-5,2,2,10,6,36,-15,0,-15,13,5,-37,5,-8,-17,-59,-7,-7,7,-25,-15,-11,-48,-5,20,53,-30,-11,12,-12,29,29,-5,1,16,-37,5,-9,-14,27,55,4,0,23,12,17,-6,6,-6,-15,-3,-63,25,-11),
	(2,-13,12,11,-36,-9,0,1,10,20,27,-25,-9,-34,-21,30,-34,43,11,-1,9,65,-13,25,-11,2,36,-24,-52,25,-3,-17,26,-13,-5,-26,-11,-21,8,7,1,-47,-23,-34,26,-30,-2,-45,23,12,14,28,14,-53,2,33,-6,17,-2,-14,5,-5,-17,-4,-11,-10,25,-7,-1,11,0,24,36,-96,-42,-25,-14,14,-7,27,-17,14,0,-9,20,-7,6,-38,-25,-24,-4,-6,10,14,-28,-44,-33,0,-7,4,-24,0,10,18,33,14,-12,4,-9,-20,18,-11,13,13,62,1,-14,13,31,7,-13,-10,-28,0,-12,-64,13,-13),
	(51,15,25,-47,-77,-20,-9,-11,-18,9,-14,14,-4,-15,-23,6,-35,9,-4,-16,46,52,3,16,17,-13,27,-40,-36,28,18,-29,6,-24,48,-25,40,-5,50,24,43,0,-13,-52,22,-8,-27,-24,26,-61,20,47,57,-33,-3,1,30,-12,4,-1,19,-32,-74,-31,-11,54,26,9,-35,55,-3,1,13,-45,-66,-4,25,-39,0,-1,15,3,-29,-45,36,-22,9,-32,-13,-15,22,8,53,-21,-7,-36,-12,-7,14,-8,6,5,-19,10,51,-6,5,9,-13,20,25,-4,19,0,16,-20,-30,18,42,-16,-5,51,-8,13,-25,0,2,-1),
	(10,7,32,11,-36,-23,6,28,14,8,-10,23,-12,-61,-26,8,-34,58,38,0,13,-4,-48,8,27,3,43,-32,-15,49,37,-44,-7,-13,34,-3,0,19,35,20,21,34,5,-17,44,-12,-8,23,52,-45,14,32,15,-16,-3,5,56,-15,-18,9,37,-1,-15,-17,-43,56,19,7,-22,23,0,6,13,-33,-24,17,25,-31,-23,14,3,24,-52,-29,43,-68,-10,1,3,-23,17,12,13,-44,-28,-1,5,-8,36,-2,11,-6,-40,44,61,16,-3,1,-33,-20,9,-16,45,8,52,-70,-35,11,25,0,-20,-2,-15,-13,-39,-25,32,26),
	(-11,-53,-24,13,-57,-2,-13,-4,18,-56,-4,12,31,-28,1,-44,-39,47,41,-22,27,-40,-46,-18,25,-2,36,-29,0,-13,26,-27,-7,-24,56,-1,-15,33,28,7,30,53,5,-37,41,-11,11,-10,61,0,-24,7,7,6,-33,32,4,-16,-21,-14,17,17,-26,-17,-24,4,-9,-5,25,12,-11,29,4,-21,0,5,20,-30,-6,19,-19,17,-22,0,16,-38,24,3,-28,-12,-18,-13,16,-40,22,-18,-18,-1,0,3,0,9,-48,-9,31,-3,-6,22,-4,-21,7,-18,1,26,34,-34,-1,-27,-6,-27,5,6,-3,-51,-2,-8,32,14),
	(-40,-23,28,-23,5,-24,3,-1,-11,-10,-21,-4,5,32,12,11,-46,-20,41,-7,44,-17,-1,-6,16,-29,-24,3,2,-1,-28,11,-15,4,9,-20,10,-11,-23,4,31,37,41,0,-4,-12,0,-26,42,-15,-10,-15,30,16,17,13,-26,-6,42,-3,-12,11,16,-31,11,33,0,-18,51,-3,-7,15,15,-23,-16,-14,-29,-25,35,-4,-37,-22,3,17,-39,37,15,0,-44,-19,-11,-10,8,-18,15,-11,-8,-9,12,50,-28,-29,0,-13,-27,-24,-8,16,-3,-16,-3,-7,-31,-20,8,-9,-29,16,-31,9,17,-42,8,-42,29,-30,22,36),
	(5,-14,18,-20,4,-21,9,4,22,20,3,3,21,18,4,-6,0,-4,22,30,30,-16,-12,-1,12,-11,-18,-8,0,2,8,-6,-9,-16,-8,-20,30,-12,-14,8,3,8,22,-8,-10,24,-1,11,9,7,-14,-18,19,3,29,7,2,28,22,-17,15,-6,9,-21,6,15,8,-5,-7,-9,-1,-3,9,18,1,-4,0,9,15,15,-20,-2,-20,-16,-6,29,20,11,6,-10,23,6,36,-4,30,-8,-4,-2,-3,4,-21,11,-17,-9,-2,-18,11,4,-19,20,19,0,-10,1,21,11,-18,-3,-19,21,10,5,26,25,8,8,-1,-7),
	(24,7,3,-17,30,7,-30,-48,-3,-7,6,-12,-7,10,14,-15,-11,2,-7,-5,28,19,25,-13,3,10,4,-2,-11,9,-7,29,0,2,3,-26,-9,14,12,-2,6,9,-9,14,-21,8,14,-18,-9,-10,8,13,-11,11,-9,-11,3,22,11,-9,-10,-3,6,-6,0,20,-9,-21,-6,6,-26,23,-8,0,-9,-21,-11,-20,9,9,-3,-18,0,18,0,0,23,6,-25,-8,-5,-9,5,12,-5,-15,9,-10,14,9,-4,-24,-15,0,-4,-19,-19,15,-13,-3,-8,11,6,23,-20,-12,-13,24,3,19,5,-8,4,3,23,0,15,-12),
	(-30,0,18,-32,9,-25,-9,-20,-10,34,-12,12,23,23,-6,-6,10,-1,20,13,-14,18,38,-14,-9,-14,-7,-18,2,20,-34,-18,-6,-27,-6,9,8,9,-16,12,13,-3,8,-2,-25,-4,27,-1,4,0,6,4,1,-30,8,-11,-20,27,6,1,20,9,-38,12,-17,36,24,-4,21,8,-17,17,-30,19,-41,-24,0,-26,-7,27,-5,-38,-27,24,-21,21,26,7,-20,19,-14,-10,-19,4,-1,-32,-7,-10,-11,-4,-5,-22,-11,26,1,0,0,28,-9,31,3,-13,-1,13,15,-19,-24,31,-30,-19,22,12,14,-12,33,-24,9,-1),
	(-37,11,15,7,-14,-12,0,-10,9,16,8,-6,0,15,0,17,10,1,12,6,-7,14,5,2,-20,-16,0,6,28,-11,-29,7,16,-19,-12,-4,-14,28,-10,-5,-15,-30,23,5,-10,12,25,-54,15,24,11,15,16,18,41,6,-8,7,-1,6,6,-28,-17,-11,-1,-31,-20,11,11,-22,15,35,0,39,10,-14,-10,26,0,26,-41,5,4,24,9,4,-10,3,7,13,-30,-50,-9,9,-12,-24,-11,-5,5,8,2,-42,-21,-17,-11,18,2,-1,-2,-33,-14,18,-10,23,38,11,17,8,-34,21,7,-33,19,13,-26,-44,4,3),
	(-19,-6,17,-19,-13,-9,-18,20,0,-13,10,35,-21,-11,6,-3,-40,30,10,-30,-4,51,-26,3,8,-1,28,-18,22,-7,-24,4,-25,-22,-8,7,3,37,7,10,38,3,39,13,-13,-10,15,-28,19,11,-4,-11,5,30,-9,-11,-29,5,-4,-2,7,-33,-24,-2,-3,5,-5,-5,14,3,-9,13,2,20,1,-19,-16,-22,-10,-36,5,6,-28,-1,-6,-1,0,7,-48,13,-4,-30,36,-14,-12,-16,-47,0,-20,10,-17,-9,-13,11,18,-12,8,-3,0,5,10,-9,23,15,24,10,-18,33,-24,-12,0,-9,-10,43,-31,-37,-20,-24),
	(-45,-7,-5,-11,5,3,22,32,26,-11,44,-7,6,-22,0,4,-18,-6,-10,5,7,11,14,-10,-18,22,-8,20,-11,-22,10,7,30,-58,-6,7,5,-5,-4,-20,-5,-28,46,10,14,-8,7,1,-13,5,-13,4,-7,42,19,21,-33,4,-7,7,-30,-29,8,-15,-43,33,-25,0,28,-7,8,-15,5,6,-12,13,4,-26,12,-29,-31,15,-27,-40,6,17,12,-7,-12,-19,-48,-6,5,-28,3,-2,-7,23,-39,37,-8,-15,-25,-13,-28,25,21,15,-6,-10,2,54,-10,10,6,-14,-12,30,-37,-6,17,-11,0,28,-7,3,0,10),
	(-39,30,-3,-20,-24,-28,37,-3,11,-23,42,7,-10,-16,15,-25,-42,0,-8,2,0,20,-19,-38,0,-5,-16,13,-26,-16,-13,-9,-4,-30,-17,-2,1,12,-43,-15,21,-8,34,16,-7,-20,-15,-28,-8,18,-39,-15,26,42,19,29,-31,25,8,0,-9,-58,-9,9,-93,-1,-39,-3,33,-8,19,3,1,30,9,17,-3,3,15,-17,-14,8,-18,-52,-14,-19,-10,-16,0,-14,-36,4,25,9,10,-27,-50,39,-14,11,-1,-12,-47,-2,-20,23,5,13,-2,-14,37,25,-18,7,46,-24,18,34,-41,0,16,-21,4,49,-13,24,-7,-12),
	(-54,27,-1,-8,-8,-12,28,-37,17,-35,61,21,-5,-27,34,-28,-34,-14,25,-44,19,-14,-19,-36,-19,2,16,-8,-1,-12,-4,21,-8,-39,16,-7,-1,-5,4,-13,15,-34,45,13,7,3,34,-4,-5,-1,-33,-4,12,44,-17,-4,0,13,31,1,17,-60,-34,12,-23,16,-30,-9,23,22,6,7,-22,16,8,14,-4,0,-3,-38,13,-4,-23,-19,0,-8,3,-26,-7,-52,-22,-3,10,-3,19,-24,-32,16,21,20,8,20,-2,6,-46,25,0,4,2,-13,1,32,-2,1,4,-28,-14,14,-27,0,-9,-24,-5,9,-14,42,-4,10),
	(-31,5,18,-16,42,-2,12,0,-21,-30,26,21,22,11,-1,6,-27,0,4,-11,-8,14,17,-63,-7,-18,18,-17,-15,-29,4,17,-11,4,14,13,4,-19,10,-9,24,-6,13,-12,-3,-38,0,-7,16,4,0,-11,17,41,1,2,-12,2,25,-10,-20,-73,-35,-10,-11,15,-42,16,38,-1,-7,-9,-34,-9,-3,13,19,-1,21,-28,0,19,-4,-2,-17,1,9,-22,8,-49,-9,-2,34,-5,6,3,-23,8,-14,11,-7,49,-16,-7,-35,-15,14,8,18,10,8,7,0,5,30,-13,-19,9,16,-5,17,-24,5,26,-14,30,10,6),
	(-10,47,35,-14,48,3,6,-27,-16,-5,32,26,12,-10,-7,-19,-35,-22,-1,-21,30,7,17,-43,20,-11,-2,-25,-11,-34,-10,1,-22,5,18,-9,-7,-7,9,-8,43,12,27,4,15,-52,-13,-2,20,4,2,5,25,30,3,0,-12,6,-3,4,0,-99,-64,-11,-3,2,-50,11,48,-3,-11,15,-30,15,-16,-11,13,-24,-2,-7,10,3,-23,16,-11,3,22,-12,-13,-60,-7,23,59,-30,35,23,-34,21,-39,29,-17,62,-7,15,-10,6,-7,-1,5,20,13,15,-7,-9,8,13,3,13,9,-7,21,-1,-23,16,-36,9,1,12),
	(35,48,21,-11,-2,-24,-4,2,-14,8,61,31,22,20,-17,9,-48,-24,11,-19,21,43,-24,6,36,5,35,-21,-10,-41,20,12,-27,-3,-7,8,12,-23,-5,26,26,-9,9,-9,-3,-45,-13,18,6,-8,-9,11,-6,35,-5,21,22,-15,17,6,8,-115,-93,0,24,25,-72,0,17,27,5,-4,-22,-2,10,-25,19,-14,-17,-1,8,10,1,-2,-17,-6,12,-27,15,-54,14,24,11,-6,-1,-7,-7,0,-32,0,-25,43,22,22,-3,-11,-8,-16,-13,7,6,5,22,11,1,0,-17,24,-8,-11,0,6,8,46,-41,27,-5,3),
	(10,3,22,-27,-45,-1,-20,-4,-11,42,43,32,32,-11,-12,-18,-34,-5,-10,-29,31,24,-14,12,34,11,15,-10,-18,-26,14,-13,-4,25,12,-12,-13,-13,5,-3,46,-3,9,-10,8,-2,-10,9,33,-39,-16,3,8,19,-12,29,9,2,20,-2,27,-118,-75,2,6,-2,-41,0,27,25,7,3,3,3,17,-31,28,-12,-9,-18,-4,6,12,-10,4,0,10,-6,15,-23,26,-5,-22,0,13,1,25,-1,-36,14,-9,13,14,8,27,-12,5,-12,-17,2,14,-4,-19,14,-2,2,5,9,3,5,-17,42,-15,23,-11,3,4,23),
	(35,0,31,-15,-49,15,-20,12,-13,44,40,-13,-13,-15,-11,-17,-31,-24,2,-40,40,12,-10,33,7,17,9,-15,-53,-18,-3,-20,6,16,17,1,-7,15,29,13,22,10,-18,-15,35,-5,-35,0,0,-53,-9,16,4,25,-4,-2,20,-1,12,-7,10,-98,-57,-15,12,-8,33,5,-7,46,18,4,-10,-12,-11,-26,13,-13,15,5,30,13,9,-77,14,19,27,-4,-7,-6,28,-9,-8,-6,-20,5,18,-5,-3,-18,-8,-22,30,-9,41,-7,13,-23,-22,13,22,-28,-12,2,-19,19,-21,41,32,-14,-9,42,0,54,-5,5,-18,-4),
	(21,-30,-8,-36,-63,-17,-14,20,24,70,17,4,6,16,-59,-5,-54,-34,16,-10,83,-15,-32,37,8,-5,-43,-6,-24,21,-16,16,-35,24,21,-33,-2,13,-32,23,44,36,20,28,10,23,-16,-39,8,-20,14,-7,-5,19,-2,12,6,18,35,-19,6,-143,-47,-34,9,-7,36,8,10,8,23,0,33,30,10,-17,-28,-20,-14,-1,-9,-15,-8,-115,18,56,-1,-1,-10,40,12,-8,0,18,8,-1,35,-19,47,-29,-7,-98,18,-19,33,-11,-7,-17,-33,-28,35,-17,-5,15,-19,-22,-19,40,-1,1,-6,22,9,36,24,-27,-29,-13),
	(-24,-49,-14,-19,0,-3,-7,1,29,-6,8,-25,14,3,-43,-19,-57,7,30,8,82,-7,-70,12,-4,16,-68,-6,-5,0,-14,-25,-1,0,39,2,10,33,-44,14,18,4,13,8,-22,22,3,-74,-17,32,21,-7,-3,14,7,6,-32,7,31,-19,17,-107,-22,-36,77,8,36,-20,-4,0,-5,0,43,51,18,10,-3,-42,14,0,-1,-28,-47,-52,16,23,-27,-8,2,58,-7,0,42,31,-6,-40,54,-9,56,-28,-6,-76,4,-1,52,2,26,-24,-58,-13,30,-38,-18,25,-31,-18,-12,25,-11,-1,-39,-16,21,-25,7,-35,-23,7),
	(-31,-17,8,-12,78,-8,-40,-1,32,-36,6,-21,15,72,3,-24,-14,-27,13,0,50,8,-62,26,-9,10,-30,-17,41,6,2,-3,-36,-31,47,19,0,12,-18,6,-7,16,22,24,-6,42,13,-53,3,-2,4,-6,9,16,14,-7,-35,9,-1,-17,22,-13,-14,-7,36,-16,38,-45,-26,-31,-5,7,49,55,-20,-1,-11,-20,10,-25,-14,-12,-36,27,-7,25,-22,-2,-1,39,-45,-10,59,31,18,-46,41,6,5,-79,-19,-28,-29,9,26,8,36,-41,-12,-27,10,-1,-4,-2,-51,-23,-17,28,7,-6,-46,-20,-1,-28,29,-64,-33,1),
	(-63,7,17,18,66,-34,-30,-16,22,-29,-33,-14,7,50,-15,-6,25,11,0,-14,65,12,20,-21,17,3,11,-4,47,-4,-20,-6,-4,-51,4,23,-19,12,-27,14,-39,-5,20,41,-30,11,-12,-23,13,38,-10,-24,-16,-5,8,-11,-21,40,-1,5,25,48,13,8,24,-5,6,-9,-5,4,0,5,73,50,-22,5,1,-14,-15,14,-19,-2,-3,33,-6,0,-15,-6,-25,0,-46,-9,75,-9,18,-21,19,15,-4,-87,-17,-17,-8,2,7,16,3,-31,43,-3,-6,10,-36,-1,-6,-5,-22,19,5,8,-55,-8,-13,-2,29,-29,-39,-4),
	(-71,7,14,-7,45,-15,-2,5,34,0,-19,-20,13,18,-18,-17,59,0,10,19,21,0,58,4,15,6,11,0,45,-30,-15,15,-9,-64,-2,24,1,10,-7,9,-14,-36,32,26,20,-1,-9,-22,3,14,29,14,21,-23,7,-10,-38,33,10,11,-1,40,37,0,-10,-20,28,-20,-6,41,0,-12,12,51,-13,-13,-22,-1,-10,10,6,16,-2,32,-6,17,-43,-25,-8,-25,-37,-12,69,-14,25,-15,11,-31,-21,1,5,-38,-23,-12,-9,4,27,-7,29,17,0,6,-5,-9,-21,-46,-14,17,2,9,-41,-20,-28,-5,-12,-15,-34,18),
	(-78,-29,18,13,-30,1,-7,31,2,15,19,-7,-1,19,12,6,38,-14,-3,18,13,-12,60,-10,14,-12,17,33,26,-17,1,7,17,-63,-16,28,-29,-16,16,-13,-6,-34,-9,18,4,-23,8,-37,23,28,1,9,1,-22,7,-4,-15,18,36,-19,-4,-19,5,8,-12,0,21,-18,-21,61,7,-4,9,5,2,-22,-2,8,9,13,-1,3,2,12,12,9,-25,-22,-24,-46,-28,4,61,-31,37,-3,-31,-8,0,32,-2,-37,-3,3,32,-5,26,-7,11,14,11,9,8,12,-3,0,13,-2,18,15,-41,-12,-4,28,9,-10,-33,12),
	(-40,-23,14,16,-17,23,0,14,25,-4,7,-23,21,36,17,1,21,-17,18,15,40,3,27,10,1,-13,18,24,-8,-39,11,14,0,-81,-18,34,1,24,7,16,-16,-16,-35,14,-6,-19,-19,-6,27,14,4,-7,30,-32,2,12,-40,22,23,-17,-15,-4,10,33,-22,-19,-9,-10,-35,28,24,-13,11,3,-36,-4,11,18,28,5,-27,10,7,14,20,21,-51,-28,-24,-51,-31,-20,74,-23,12,-7,-78,-16,3,59,5,7,-11,32,20,35,31,-3,14,-10,22,1,-12,-5,9,0,3,17,-6,-19,-72,-6,-36,5,12,-7,-29,20),
	(-41,10,-5,17,-53,-15,21,-11,-8,1,32,-20,-18,-4,-1,-1,-26,-1,-9,4,22,54,19,10,-1,-15,32,29,-32,-15,-4,12,4,-62,2,11,-11,21,16,0,-23,-32,-53,-42,-12,-25,-11,-18,37,17,-3,-5,38,0,-18,6,-27,24,15,-19,17,3,25,9,-51,-5,25,-18,-5,33,-5,21,39,-29,-37,-10,-7,29,5,16,-15,-4,17,13,-3,4,-10,-44,-37,-20,-20,16,76,1,-4,-9,-31,-20,-1,67,1,-25,12,7,24,29,21,-10,1,-4,3,-5,-24,19,47,41,0,-3,-3,-15,-53,-22,-32,21,-17,-32,-14,-8),
	(-45,-31,19,12,-44,7,15,-29,-18,27,1,6,-23,0,17,-12,-11,8,2,-5,17,54,-6,13,12,-21,17,-1,-58,16,10,-2,-14,-102,4,-19,-19,-19,29,14,-31,-37,-31,-71,8,-6,4,-33,35,-4,-5,1,6,-39,-34,39,-42,0,21,-9,14,-23,13,-3,-44,6,39,-14,-29,19,-1,42,3,-48,-27,-27,-13,27,27,33,-13,-11,4,-13,17,-16,-3,-40,-2,-64,6,-4,46,11,-30,-18,-39,16,-19,60,-8,-10,4,15,35,10,-6,-9,18,3,-2,25,-6,4,26,19,-26,20,9,17,-43,28,9,36,-17,-42,-13,6),
	(-53,-33,1,30,-10,-6,10,-17,-10,26,-13,-35,3,-10,14,4,-17,14,11,28,33,62,-1,7,-3,-6,-2,-4,-23,12,-3,35,10,-85,-20,-40,-16,-16,33,-11,-6,-5,-18,-46,-10,-26,11,-39,25,12,42,6,23,-5,-6,22,-24,22,12,-5,27,-10,-22,-14,-23,11,53,-36,-25,-7,-21,26,41,-69,-26,-1,-31,9,4,46,15,-2,5,-6,18,-27,-12,-72,-36,-15,-9,1,12,6,-28,-3,-26,-6,8,29,-32,4,18,0,-3,38,0,5,4,-15,17,18,0,15,47,38,0,19,16,11,-39,-17,4,27,-8,-54,-6,2),
	(-24,1,-24,3,-10,-28,3,18,17,38,14,-3,-28,-2,-6,12,-51,16,4,-6,8,25,0,24,-5,15,34,8,-27,8,-4,1,11,-33,-13,-19,-27,-23,24,-20,-15,5,-28,-52,4,-19,-6,-38,-6,-14,19,32,16,-21,-6,6,19,13,17,15,29,0,-44,8,-43,-23,40,-9,-2,-6,5,-3,56,-75,-1,0,-10,-14,-3,11,6,2,-8,-51,29,-6,-22,-34,-17,-26,-36,40,22,19,-20,4,-5,14,29,4,-20,-1,45,28,20,43,11,13,-9,-33,29,3,12,-7,7,24,14,11,31,-16,-71,-2,-38,6,-31,-41,-16,14),
	(-49,5,10,-34,-70,-5,-1,-5,-26,-1,-10,0,13,17,-13,0,-43,2,-4,-8,53,9,-1,2,37,-9,35,-41,-26,44,0,-28,17,-37,11,-34,20,-12,47,-4,15,12,-38,-42,4,-19,-1,13,31,-46,-17,41,28,-32,-4,-13,21,-44,-25,0,6,-15,-70,-25,-6,54,52,10,-35,11,-19,-5,32,-62,-16,-19,49,-25,-11,-13,17,9,-35,-34,-4,-4,-26,-3,-26,-42,-20,15,84,2,-31,-9,2,7,31,-8,-1,5,-33,1,48,8,-22,23,-15,-13,15,2,16,-58,-4,-18,-26,-12,72,-16,-50,23,-2,15,-43,0,5,-3),
	(13,13,43,3,-52,-49,-7,-2,-3,-27,-5,-6,20,29,-4,-8,-24,13,5,25,22,-15,-18,-15,10,-26,33,-39,-18,25,31,5,8,1,10,-33,4,5,35,5,8,23,-6,-11,22,1,-22,3,44,-38,-18,14,-7,4,0,-12,46,-11,-36,-10,9,18,-13,-22,-23,29,42,-32,-6,20,-46,-3,51,-2,-15,20,13,-29,-22,-29,23,33,-32,-18,13,-26,19,18,-35,4,0,-32,44,-62,-22,-26,30,-1,3,0,15,-24,-47,-25,24,-32,-2,11,10,-12,18,3,-22,-25,1,-60,-43,3,51,15,-5,12,-1,-47,-37,-3,35,52),
	(-12,-37,30,10,-23,-3,-23,-26,6,-54,0,23,8,-15,-21,-11,-44,12,26,-1,44,-26,-34,-35,19,0,27,-25,1,12,19,-6,20,7,54,-24,7,25,12,9,27,39,28,6,17,-30,9,14,40,-14,5,41,3,36,-2,-4,11,-26,-42,-19,25,0,8,-30,16,17,31,-3,29,36,-22,12,37,-10,-16,10,8,-11,-24,-30,-6,-9,-27,-13,14,-6,32,-6,-51,16,-23,-15,40,-15,-7,-41,7,28,17,-17,22,-19,-8,-2,29,-23,-11,-14,-21,-32,9,0,3,7,-3,-27,-34,10,-4,25,7,11,2,-26,-11,22,46,25),
	(-12,21,-1,-13,27,-18,2,-5,17,-24,2,4,33,18,0,-4,-11,7,9,-12,32,10,15,20,-14,-6,1,-10,-5,-20,-7,11,-8,2,-7,9,16,-25,-40,26,22,20,20,-6,-36,6,36,4,33,3,-1,-2,15,16,-19,10,-2,-17,42,16,-28,22,14,-28,25,23,-29,-40,52,-13,-8,10,10,-10,-11,-5,1,4,22,18,-49,-33,-27,18,4,22,16,-6,-37,17,-3,-14,-34,-9,24,5,-1,-29,0,57,-25,-23,-9,3,0,8,9,8,16,-25,21,-10,2,-9,14,13,-21,0,3,23,-9,-23,30,-3,-9,-30,27,27),
	(-13,22,12,2,-16,-26,15,-19,3,14,-35,8,4,22,7,3,12,-9,-2,4,17,19,-1,7,38,-16,9,-17,0,4,-7,19,-11,2,22,-13,10,-18,-5,34,24,21,8,-21,-31,0,24,-21,17,21,-5,-5,-5,3,-6,17,0,7,14,-4,-7,-18,-3,-15,-27,7,-9,-11,27,31,-4,8,11,8,-17,-4,-12,-28,29,-7,6,-9,-8,6,-5,0,33,-5,0,9,1,-25,19,2,3,0,10,-21,14,18,13,-21,10,-39,-7,-8,14,39,10,31,26,-18,-21,22,2,5,-30,17,-11,-18,26,-20,-15,16,27,9,8,-7),
	(-36,2,-10,-17,3,-19,-14,-39,-24,29,9,-6,0,2,-3,-15,17,13,26,30,11,30,48,34,4,-26,22,-21,7,-7,-11,26,2,11,10,-25,-3,9,-16,7,5,0,21,25,-29,19,24,9,-2,3,20,16,35,12,-14,-37,-27,5,28,-11,20,5,36,-17,-3,22,22,-4,46,39,-22,12,-5,3,-1,3,-15,-2,2,9,9,-21,-25,14,-27,18,21,8,-26,21,-8,-3,18,37,-1,0,-37,-48,-8,-12,1,-10,-1,-1,3,45,-24,-7,-10,29,-13,-22,-23,15,-35,23,-28,31,-13,12,19,18,-24,7,25,-21,12,-48),
	(4,-16,8,-5,6,-27,-14,-29,20,28,-31,-11,7,16,41,-20,12,-1,20,-7,34,38,-12,-31,22,-18,-23,1,20,21,-40,31,-21,8,5,-34,0,7,-28,47,21,11,14,-46,-6,-17,-2,-26,39,18,-2,2,32,-12,-8,19,-9,28,2,15,13,-21,-47,-20,12,31,18,-7,-2,20,-24,-4,3,12,-18,-32,-31,-15,33,27,-35,-14,-15,34,-30,11,32,1,-14,11,-8,-14,24,-12,28,6,-20,-7,5,16,-7,-30,10,-39,-2,-19,-4,25,-11,11,27,-19,-16,32,27,17,0,-4,-34,16,10,-5,7,28,20,-38,0,-29),
	(-12,-12,-6,-8,0,-18,13,55,39,9,4,5,7,-5,0,-11,-2,18,-5,30,4,0,-15,-3,-8,-2,-21,14,-1,-2,-35,45,-5,0,-6,-11,2,5,-2,0,14,-22,38,-11,-10,4,10,-30,33,47,3,-23,16,-3,8,-1,-37,13,-3,-12,11,-19,-33,-5,-27,1,17,-14,-10,17,30,38,-5,21,3,-39,-28,-33,-22,22,-25,-15,-15,12,11,0,-15,-7,-21,49,-16,-16,-1,22,13,-34,-8,23,42,14,7,-28,-32,-6,-15,35,5,-4,-19,0,8,9,0,58,17,-18,1,6,-55,12,-16,-25,-33,15,3,-8,-15,-12),
	(-13,-12,-34,-15,-28,7,-4,38,17,-23,51,16,-4,-8,-8,-28,-22,9,17,-21,14,23,-24,-6,-4,-8,-4,-3,-4,-16,-15,30,-8,-23,15,7,-24,23,-33,-22,38,11,30,-2,-1,-17,16,-23,6,10,-56,-28,20,42,5,7,-3,-1,10,-12,1,-75,-26,-32,-24,-15,5,-12,-23,-7,0,8,-2,17,56,-27,-11,13,5,-36,-41,-18,-28,-10,27,-30,15,2,-46,-22,-37,-22,13,-9,-13,-40,-58,20,7,37,-19,-18,-10,33,8,-1,13,10,-20,-18,0,11,14,35,34,2,17,7,-60,-3,33,-21,-3,40,-35,-44,-49,-10),
	(0,15,12,4,-19,-7,10,48,-23,-47,53,19,27,-33,16,-38,-11,0,-22,-6,-7,25,-17,-33,5,6,25,-15,-10,-14,18,-5,10,-39,-22,2,8,-12,1,-8,15,-6,25,0,-4,-41,10,-13,5,9,-60,-16,10,23,0,36,-31,-53,-15,-14,-5,-57,-40,-4,-27,5,-29,-11,21,-32,7,-15,-6,-4,20,-13,12,-1,18,-24,6,42,-5,-26,-9,-37,8,-15,-45,-27,-26,-28,6,-47,27,-24,-8,52,-26,34,13,0,-39,10,-3,3,27,-2,-21,-25,43,23,13,1,21,-19,2,4,-40,-22,29,2,0,60,-26,-9,-13,20),
	(-46,20,10,-5,-18,-8,11,-21,-18,-23,48,46,1,-12,-11,5,-53,-1,14,-19,-2,34,21,-44,13,-11,5,-16,-5,-16,0,-1,-6,-25,19,-17,22,-23,-4,-10,3,-18,20,8,-1,-34,21,-40,-14,-18,-47,-7,12,24,0,28,-31,-11,10,-18,-29,-60,-48,28,-62,29,-31,37,2,-20,0,-44,-44,-6,11,2,13,6,-18,-1,8,20,-12,-28,-30,-42,18,-45,-20,-43,-52,3,0,-29,43,-17,-3,14,-38,42,9,21,-4,20,-24,0,19,-12,-4,6,8,38,0,-21,12,-5,22,19,-14,-14,15,7,17,25,-18,31,12,17),
	(-32,24,15,14,-1,19,18,-48,-23,-4,64,0,-3,-23,1,-16,-17,6,20,-56,22,-5,9,-41,12,-5,6,-35,-6,-9,-16,12,-25,-27,15,-9,-7,-31,2,1,32,1,-2,-15,-15,-5,21,-16,7,-4,-22,-11,45,22,-33,24,0,-4,21,-14,-5,-106,-54,16,-18,11,-31,-1,-6,4,8,-8,-10,3,2,-2,19,9,22,-12,-6,1,-15,-17,-29,-21,27,-26,-4,-31,-35,26,1,-9,48,-12,13,9,-8,52,3,15,-17,-1,-34,28,29,31,-23,-15,14,0,-20,7,-13,-14,2,24,5,-17,-8,11,7,42,-14,42,6,-5),
	(-2,15,22,8,19,-24,16,-10,-27,-3,37,15,-18,20,29,-32,-24,2,9,-22,26,19,0,-36,4,-14,1,-11,-15,-13,-9,8,3,-12,5,-19,4,-13,-3,-21,29,19,-11,-16,25,-34,14,-20,0,21,-13,-9,12,17,-5,27,9,-10,29,-22,14,-100,-58,29,9,27,-37,19,-27,-3,-16,-9,0,-14,-9,7,26,-7,13,-30,9,28,-4,1,-22,-5,17,-25,17,-45,-36,31,49,-13,36,34,-5,44,-30,42,3,42,26,-14,-24,-10,25,0,12,12,16,1,12,-25,25,26,-5,17,16,-33,3,-9,0,43,-28,12,-6,-2),
	(-1,55,22,-10,22,9,10,-17,-30,22,30,27,-19,0,2,-45,-25,-25,6,-32,14,23,6,-38,15,12,14,-3,-27,-53,0,1,-25,1,10,-22,-5,-6,-9,6,10,15,-10,-18,10,-9,23,5,13,17,-16,13,30,-18,-8,11,0,-20,21,-23,-2,-88,-75,0,-7,36,-30,11,-11,2,3,-16,-16,-3,-26,-28,25,-14,4,16,-19,-5,0,12,-16,-15,42,0,17,-16,-2,-4,32,9,28,25,20,23,-55,16,24,68,-5,-10,-10,0,20,4,-7,17,20,-28,13,-14,17,-10,2,-22,17,-19,8,-22,-21,45,-27,14,8,17),
	(-7,33,18,-20,-17,-5,-12,-23,5,47,2,9,-16,-13,-1,-47,-38,-33,7,-36,18,36,-4,-5,-2,-30,29,-37,-10,-31,-7,3,-14,22,8,-18,13,-30,9,10,23,1,-12,0,1,-6,2,7,36,-8,-26,-15,10,-1,-18,2,2,-7,33,-9,2,-77,-68,10,26,-3,-44,8,-62,28,-13,-7,-9,1,16,-34,-12,-35,35,6,6,6,14,-21,-6,0,22,-11,29,7,20,-9,13,-10,22,6,36,5,-43,19,-13,39,13,-24,-19,-31,16,9,-30,0,29,-13,-16,-9,4,8,-7,11,1,-38,-1,-4,5,68,1,8,-16,18),
	(24,-22,17,6,-38,-14,-24,35,-2,82,-7,39,-24,0,30,-38,-38,-16,-1,-36,39,16,4,-1,31,-21,32,-13,-30,0,-7,-29,9,0,10,-13,7,-23,8,20,23,13,7,4,34,-2,-15,16,28,-10,-5,0,21,-10,22,22,10,-14,4,8,15,-68,-19,2,3,9,-31,-20,-58,7,-19,-38,6,-9,-15,-4,-11,-11,23,11,14,8,-7,-58,-21,30,39,-11,16,27,6,0,16,2,3,0,45,-1,-27,-32,-12,11,-9,8,4,-23,-3,-8,-30,-1,4,-38,17,13,0,2,-10,9,-12,-9,-31,2,13,86,-1,6,-32,0),
	(0,-29,1,-35,-55,-18,6,19,-8,71,-25,0,-44,-4,-26,-38,-17,-60,-40,-8,8,8,-10,32,-2,21,43,-16,-25,8,12,-22,-11,18,12,23,3,-7,-9,-4,-7,19,-6,4,36,47,-21,1,0,13,20,22,-25,-3,-1,28,23,-1,18,8,22,-58,-20,-16,14,25,12,-10,-97,44,0,-12,-11,1,27,32,16,-48,8,17,4,8,12,-117,-17,50,10,-4,25,15,6,22,13,10,22,-16,27,-6,28,-9,-32,8,-3,7,35,-10,5,0,-35,30,9,-38,25,36,-42,-18,-8,9,25,-16,-39,35,-2,57,42,-11,-43,6),
	(-21,-46,11,-33,-13,-21,-23,19,-9,39,-51,-15,3,-6,-50,-47,-25,-28,-15,-11,58,-9,-54,21,19,5,-20,-54,0,35,-5,3,-12,11,3,5,-6,22,-31,7,9,30,20,19,-1,36,22,-35,41,31,12,-28,2,60,-24,-1,15,19,19,6,47,-78,-19,-15,35,-5,11,16,-81,-13,22,-24,38,13,22,44,-12,-53,10,-10,14,-31,-41,-96,10,27,0,13,-6,51,-7,34,-1,22,-5,-6,34,-14,33,-9,-34,-26,8,28,47,10,20,-27,-33,6,24,-50,19,32,-59,0,13,12,11,-8,-48,25,5,7,43,6,-36,21),
	(-22,-35,-16,9,12,-1,-31,-14,0,-45,-35,-7,5,46,-42,-42,-15,-18,-13,-5,75,23,-59,51,-22,31,-49,-50,30,21,2,14,-12,-10,27,38,-16,20,-33,-9,-33,31,33,11,-1,23,28,-37,25,40,25,-17,17,48,1,-2,34,21,-3,7,30,-43,-28,-28,74,0,42,1,-39,-58,3,-9,53,36,33,28,5,-52,1,-18,2,-38,-49,-1,24,17,-27,-4,-37,27,-16,-9,41,29,-1,5,46,-16,20,-32,-27,-52,32,28,30,-11,37,-34,-29,-28,36,-51,7,21,-52,-17,16,-11,-7,-16,-56,-22,27,-60,20,-13,-28,4),
	(-46,-34,5,-15,53,-9,-31,-34,31,-57,-21,-19,-8,29,-9,-38,5,3,1,-46,16,9,-29,-3,13,5,-21,-12,50,-14,25,11,-8,-28,5,35,-21,28,-21,0,-53,38,13,29,12,22,18,-30,17,13,3,-27,-18,-9,-2,24,20,6,0,4,23,13,-4,14,50,-3,31,-24,-17,-32,-2,0,43,46,37,1,0,-26,18,-8,-35,-1,-36,52,-2,0,-28,7,-28,25,-23,-3,50,-4,16,-1,-10,-25,25,-34,-47,-32,3,-16,0,-26,17,-34,3,-14,0,-25,-2,17,-18,-34,-23,-2,-2,-8,-62,-6,46,-33,13,-47,-28,11),
	(-49,3,31,-10,18,-19,-30,-7,22,-12,-17,-22,8,29,14,-30,38,-28,10,-20,7,-7,18,27,13,6,-18,-5,17,-52,-10,14,-10,-38,6,17,-2,11,-8,8,-35,17,29,31,1,-12,-10,-5,10,24,17,-15,-21,4,27,-10,-3,-21,10,-17,13,27,-3,12,29,-6,11,-29,-16,-31,-6,-38,3,-5,17,5,18,-32,21,1,-28,-14,-20,19,7,16,-9,26,-26,-27,-19,-14,57,-48,37,1,-5,-2,0,-11,-11,-33,-19,7,-4,-32,7,-32,23,-26,17,-15,-10,15,-27,-43,2,-32,-7,-12,-18,-28,17,-23,26,-25,-42,26),
	(-77,0,1,-8,14,-17,2,-3,12,6,-18,-25,20,34,7,-11,32,-9,-10,14,-10,7,38,-7,12,3,-9,5,9,-44,12,27,1,-10,-24,29,-19,-7,-6,-7,-11,0,20,11,-8,8,-10,-6,21,40,-3,-13,12,-5,3,10,13,16,15,-15,13,35,26,19,34,-3,9,9,-10,1,25,7,15,43,13,2,-22,6,17,7,-4,18,11,22,13,20,-6,10,-44,-38,-13,19,65,-52,16,1,-36,7,-16,43,-22,-32,-8,9,-10,1,13,1,36,-12,11,10,-5,-6,12,-51,9,-4,31,20,-24,-27,38,30,7,-7,-26,11),
	(-67,13,-8,16,-33,-16,2,10,3,12,3,-11,6,39,-5,-29,8,-25,0,11,14,-10,30,3,-12,-14,9,27,-20,-20,-18,33,16,-16,-21,29,-3,-3,1,-14,15,0,18,17,4,-13,-3,-2,-7,20,-31,4,-7,16,20,9,-26,-8,9,-6,-14,14,7,31,25,9,25,-4,-27,43,2,18,-13,19,6,2,-10,21,-17,-19,-14,26,-22,-2,1,22,3,0,-24,-28,-24,7,77,-33,25,17,-38,15,11,32,-35,-3,-14,-7,12,13,-2,20,20,9,14,13,-28,-6,22,-14,-19,7,-1,-9,-36,-26,-13,16,8,16,-48,22),
	(-87,-33,-32,28,-49,23,28,-13,10,-5,14,0,4,26,22,-12,-4,8,3,18,0,20,25,-6,-21,16,31,39,-27,-20,-9,37,1,-31,-21,26,-18,0,-9,5,-14,-1,-18,20,-3,-29,-18,-17,-8,9,-9,28,-3,-15,-11,-1,-44,2,17,-3,-22,-9,22,9,-25,-5,0,7,-33,29,5,-16,-3,0,-21,-26,-10,14,-3,-3,6,2,22,-25,24,29,14,-6,13,-13,-34,3,37,-3,2,19,-72,4,20,41,17,-23,-12,9,-7,4,20,22,26,17,28,19,9,12,31,12,5,13,16,13,-56,1,-26,18,31,-14,-31,9),
	(-71,3,9,32,-34,-17,27,-1,10,12,-10,-25,-17,34,2,0,-33,9,-22,4,18,45,14,-7,8,14,12,41,-41,-35,-26,38,16,-28,-13,0,-11,-17,3,-23,-25,27,-16,15,-16,-10,6,-27,-27,14,13,-16,17,-4,-39,31,-13,28,38,17,-8,1,37,-5,-37,3,-12,-16,-39,-1,19,17,19,8,4,-10,-8,18,-2,-9,-28,32,-6,-24,12,13,0,-30,18,8,-22,13,46,4,0,25,-24,9,-13,45,5,-19,3,21,-14,6,9,42,24,16,0,34,-27,-1,32,29,16,-7,18,13,-78,-15,-15,19,23,-18,-39,6),
	(-72,5,-19,23,-29,-9,31,-34,-5,-15,-2,-2,-27,4,23,-16,-43,-14,0,-15,29,55,-4,-6,17,5,-20,2,-37,-13,-23,25,2,-59,-1,-23,-40,-48,-7,-49,-18,-18,-6,-26,3,-42,25,-6,-15,16,16,-6,24,3,-61,19,-12,15,19,-18,19,-16,0,0,-10,2,16,-1,-20,5,13,3,9,-16,-3,-25,7,46,0,13,4,10,8,6,-5,-7,-11,-39,0,-3,-24,0,42,16,-11,-7,-3,3,-41,29,9,0,15,-10,-8,-1,12,22,28,12,-5,32,-14,11,19,19,-19,-13,9,-32,-74,2,5,14,14,-36,-32,8),
	(-106,-21,-4,4,-32,-9,6,-14,0,-5,-19,-26,14,-30,19,-10,-13,-3,19,-6,52,55,22,34,3,9,-2,1,-21,-4,-40,33,3,-79,3,-18,-39,-70,21,-31,-24,9,0,-60,-4,-41,-10,-27,-2,-1,14,-7,1,23,-28,-3,-37,46,34,-4,2,-6,-21,-19,-39,-18,35,-1,-14,10,15,-8,30,-53,-10,-26,0,9,35,5,-19,-11,5,7,-3,-25,4,-50,-36,5,-21,-20,69,-4,18,-8,-10,28,-19,25,-8,13,15,0,-2,20,-1,17,18,-22,12,27,-39,7,22,16,-1,-18,23,-4,-79,7,-24,-2,9,-15,-25,-9),
	(-91,1,-9,-7,-4,-8,-2,3,8,29,-16,0,14,-9,10,-14,-53,26,20,-36,39,27,-2,35,20,-2,13,0,-21,10,-28,38,21,-33,-1,-37,-24,-28,4,-33,-14,9,-47,-57,-12,-33,13,-23,-4,0,-5,1,29,7,-31,0,1,-2,24,-5,11,-32,-51,-24,-33,-11,42,31,-5,10,-6,-29,27,-34,4,-17,-19,23,-14,8,-6,23,-36,-40,-5,-46,-15,-54,-15,-3,-37,-1,54,27,-5,24,0,15,-8,-50,8,19,5,-1,49,20,-4,-1,-23,-36,3,9,-2,-23,-11,13,7,-17,71,-10,-96,20,-10,-18,-17,-34,-33,13),
	(-50,16,-24,-31,-62,-4,-11,5,-1,12,-4,46,2,16,-26,29,-67,30,21,-3,39,-6,7,-5,54,-4,9,-3,-2,5,26,18,12,-22,26,-35,-29,-16,50,-46,2,19,-56,-54,-1,-55,-1,-9,8,-52,27,7,56,-7,-53,-30,27,-7,-3,-8,7,-9,-62,-43,-44,38,30,31,-30,34,23,-17,52,-57,0,-19,28,-13,-36,-12,10,21,-58,-63,8,-50,-11,-44,-41,-70,-59,1,108,18,-23,11,23,9,-15,-51,38,42,13,23,67,36,-22,2,-40,-37,18,19,24,-41,0,0,26,-18,76,-32,-49,27,-40,-19,-68,-13,8,20),
	(7,-17,2,22,-43,1,-3,27,24,-9,11,8,-22,18,-25,6,-62,40,11,5,66,-23,-30,-8,34,29,40,-21,-28,-19,41,-18,40,-11,45,-23,-10,-1,29,-8,-13,18,-42,-33,29,-41,-32,4,-6,-52,1,10,11,3,7,15,26,-9,-67,-13,12,-27,-3,-57,-51,-9,36,-4,30,18,12,11,45,-16,-17,34,52,-22,-47,-27,-18,47,-15,-39,17,-56,-35,-7,-50,-16,-53,8,27,-57,-9,-21,35,38,-23,-13,56,0,-31,23,56,5,-2,-31,-3,-43,18,10,3,-9,-24,-14,4,24,30,-8,-22,26,2,-62,-27,-34,5,16),
	(-12,-48,13,1,-42,-14,-5,-25,16,-34,14,49,-17,-28,-55,-22,-25,3,-1,8,38,-48,-25,20,31,27,44,-31,-1,15,56,-12,35,-8,64,9,-5,24,12,24,16,37,-40,-23,54,-23,-12,22,34,-4,41,64,14,46,-22,28,24,-37,-22,12,62,-49,-9,-19,-31,30,26,9,5,28,14,20,2,-18,17,-12,31,-10,-17,2,19,41,-26,-53,0,-74,-1,-1,-18,3,-21,2,38,-27,0,-33,-2,34,-16,-10,-10,14,-18,5,55,23,10,-41,-15,-63,22,11,16,12,16,-61,-9,48,46,10,-15,-7,-32,-20,-53,4,22,37),
	(-27,35,23,-6,7,-22,15,-21,33,1,16,18,17,-15,-17,-14,-5,0,13,-25,28,20,-20,-7,12,0,-28,-26,-4,17,-3,0,-9,-19,23,-20,2,-10,-33,28,14,40,-6,-3,-21,2,17,-12,9,-18,12,0,33,22,18,28,18,-2,16,9,20,7,-7,-26,6,-8,0,-13,-16,4,-5,4,22,-15,15,13,-22,8,-20,-2,-36,-2,-37,13,9,-20,-11,-16,-43,21,-17,9,18,-23,26,-1,10,6,-11,37,-28,-17,-4,1,21,-5,23,2,-3,10,9,5,-11,-28,13,-29,-7,9,-10,6,8,-19,-1,6,-21,-14,-21,9),
	(-16,8,14,-18,22,-20,5,6,-18,-7,-15,18,-15,-14,0,6,1,-4,31,-11,31,31,4,-7,10,-11,16,-23,28,17,-3,0,-7,8,-15,-20,31,-3,20,15,34,-10,0,0,-17,14,-13,18,32,-4,-18,-14,8,5,16,-2,-6,1,26,18,-4,-14,-15,13,9,3,14,-14,6,21,-34,-9,-1,-5,-20,7,-15,-6,4,-1,10,-5,3,11,2,24,27,-7,-12,14,9,-14,-14,16,21,5,-7,-23,14,-3,14,6,-1,-21,6,-21,-4,16,31,6,-3,-28,-11,21,8,-16,-31,-4,15,-3,18,-10,-16,17,20,-9,18,1),
	(-14,13,1,-17,16,5,5,-26,-15,-4,5,0,-4,22,13,-16,-1,5,27,27,-4,65,13,5,11,-16,16,-10,0,26,-10,9,-26,12,-1,-18,6,11,-6,3,0,15,-7,-3,-12,11,-6,-16,-1,7,-18,0,-6,8,19,2,-21,14,11,14,6,0,-8,-4,-16,4,2,-20,22,-4,-2,2,12,2,-11,6,4,1,-4,-5,-3,-14,-24,-4,-12,-2,32,-11,-15,13,-8,-31,7,4,-11,-1,-31,-30,24,28,-21,-3,-2,1,19,-10,-19,10,-7,-10,-4,-51,-22,10,2,4,8,-6,-22,-4,-7,-9,5,36,21,-21,-4,-11),
	(-9,-1,0,-26,18,-8,-5,-15,0,10,26,-3,28,40,10,-28,-10,-6,29,-8,37,7,0,-37,17,-25,6,2,40,7,-22,14,-28,-4,21,-20,13,-4,-15,30,42,18,27,-27,-24,-14,-3,-38,33,24,-39,-27,9,2,4,-6,-26,9,9,0,-6,-39,-26,-17,18,33,32,-2,-18,7,-34,-10,21,10,-22,-16,-31,-9,4,4,-14,-13,0,16,-34,15,24,2,-6,27,17,-45,18,22,17,9,-21,-13,-5,40,-13,-18,3,-31,17,0,-31,-11,-34,0,20,-22,-35,35,-8,-3,-25,-7,-18,-2,17,-18,17,3,23,-22,7,-9),
	(-9,9,7,-3,15,0,12,33,13,35,0,13,-4,26,-17,-24,-40,-9,-11,-29,-4,11,-28,-17,-4,-12,17,-3,-9,-21,-12,6,-3,-22,-11,-25,-8,17,-22,0,10,1,49,9,-32,-14,0,-13,11,50,-26,-12,27,16,16,13,-9,-5,30,-20,10,-58,-32,-35,-17,6,7,-21,-48,24,23,4,30,18,-11,-22,2,-32,-8,-16,-28,9,-48,0,5,-8,0,-31,-28,-2,-35,-2,23,-18,7,-6,-48,-11,26,17,-36,-16,-29,-8,-10,20,16,20,-15,-28,32,16,0,28,28,-34,-27,2,-38,16,-28,-10,8,8,-5,12,-15,3),
	(23,12,-24,26,-25,-11,-1,62,-20,-33,50,-2,-42,11,-11,-25,-35,0,-15,-44,12,21,-6,-8,19,15,-10,-14,-11,-19,16,32,-3,-10,-11,2,-13,6,-38,-17,32,32,24,29,11,-5,-1,-35,8,0,-59,-4,16,34,-20,28,-35,-9,22,12,51,-95,-42,-31,-28,-4,-1,-18,-63,-32,22,-17,19,28,10,-9,-11,-5,-28,-22,-14,17,-36,10,11,-42,42,-10,-58,-21,-43,-27,12,1,31,-31,-56,12,29,39,0,-24,14,1,9,22,11,25,-24,-24,9,32,-14,7,7,20,-4,22,-31,15,-20,-2,12,42,-37,-22,-41,23),
	(-10,7,-4,11,9,-3,12,14,-11,-2,18,7,-18,-34,12,-43,-15,-7,-23,-31,-9,35,-8,-20,14,17,0,-24,-9,7,-3,3,-2,-39,-9,-17,-22,0,-25,-11,-5,-1,38,-17,31,-30,-22,-34,26,13,-59,-14,-1,14,-41,17,-37,-35,4,13,32,-82,-33,3,-49,15,-23,-3,-42,2,33,-26,-25,8,20,-10,-11,-28,-11,-29,-13,22,-32,-43,-23,-47,46,-14,-45,5,-25,-22,8,-37,45,-17,-1,13,-29,10,3,13,5,-2,-4,4,44,6,-28,-22,27,11,4,0,3,-5,0,17,-32,-22,-25,-19,18,55,-46,-11,-39,12),
	(3,45,9,7,9,-4,31,-13,-68,28,28,18,-15,-1,-9,-50,-19,-14,-21,-35,11,16,37,-32,21,9,3,-29,-23,-9,13,0,-10,-46,-26,12,-2,-16,21,-8,32,8,-11,-33,26,-16,-15,-29,19,-18,-10,9,5,19,-46,6,-19,-38,32,-2,0,-68,-64,26,-39,36,-29,35,-29,-6,4,-32,-23,-7,9,16,-18,-15,-6,-33,6,22,-24,-32,4,-48,38,-7,-14,-16,-14,11,-1,-10,5,0,14,-24,-48,37,18,29,-17,16,-28,30,18,8,2,-30,4,30,5,3,8,1,18,10,5,-17,-19,-5,7,1,-33,37,-27,14),
	(0,11,37,6,19,9,-3,-23,-56,13,28,24,0,-11,31,-45,-20,-2,10,-56,16,14,10,-27,0,-6,8,-11,-11,-31,-4,6,-6,-29,2,-13,8,-13,-6,5,2,13,-7,-25,5,2,-22,-23,13,-21,-26,-4,24,6,-21,2,-2,-30,9,11,4,-97,-57,1,-1,14,-11,25,-71,3,10,-33,20,20,-22,15,10,-21,12,-26,-5,-4,9,-20,10,-2,18,-10,20,-12,-11,9,31,-5,20,-21,5,12,-33,22,2,15,11,27,-24,24,10,14,13,2,3,3,-3,-22,9,-18,1,28,5,-27,1,-6,-13,35,-30,8,7,-11),
	(-6,27,27,14,33,-8,-12,-35,-34,50,34,8,-33,-6,43,-47,-40,-20,16,-25,5,54,-2,-53,12,-2,-6,-9,-15,-14,-16,-14,3,-4,0,-6,-11,-32,7,-13,-3,4,-4,-16,2,3,5,-8,22,9,-33,6,-2,21,-13,15,-17,-4,14,-1,-9,-76,-43,6,-8,44,-41,18,-79,22,-28,-21,19,0,-20,22,1,-26,8,0,-14,-13,3,-4,-26,-7,31,-2,26,-12,-11,0,16,5,19,10,21,5,-29,12,29,12,-13,-3,-11,-8,8,-2,-5,4,18,18,-10,-13,-2,-4,-7,17,19,-37,-12,0,-3,42,-24,16,-2,-13),
	(7,12,41,14,15,26,26,-14,-32,87,18,22,-14,2,0,-40,-35,1,11,-28,-4,44,6,-9,-5,-6,14,-7,-8,21,6,-16,9,26,4,-8,-13,-7,-8,15,12,0,-13,7,-4,6,-20,2,25,-9,-20,10,20,-2,2,4,-16,-12,15,-14,-8,-57,-65,26,29,0,-28,24,-98,9,-22,-39,4,5,-13,6,15,-17,-3,8,-7,17,22,-60,-9,-1,19,21,11,15,-12,-6,24,23,0,20,38,15,-32,-7,28,43,-2,6,0,-11,4,-4,-25,18,12,-11,19,-12,-24,2,0,12,13,-29,-3,-37,5,37,-9,6,-9,1),
	(22,22,14,15,13,4,12,-2,-14,87,-31,41,-27,-15,8,-16,7,-15,-19,-31,-11,26,25,6,15,-27,48,-21,12,5,-2,-7,29,16,8,-8,-4,8,31,9,18,6,-24,-15,30,27,-28,0,38,-25,13,10,19,-25,18,-11,18,0,19,5,10,-31,-24,0,32,5,6,19,-68,26,-13,-36,5,-7,-17,34,15,-16,2,7,16,-4,-9,-66,-3,22,23,39,5,18,38,5,12,15,13,16,34,0,-14,-25,1,61,10,6,-32,-36,19,0,-5,28,-23,-9,5,10,-1,16,3,9,1,-20,-34,-5,-5,55,2,-16,-21,3),
	(15,-57,8,-10,-43,-2,-19,28,-4,83,-56,23,-42,-11,9,-30,8,-43,-53,-25,-30,30,-13,9,15,0,47,-31,10,15,5,-9,7,8,1,34,-7,-26,27,-6,-6,-17,-28,11,32,55,-33,44,12,-15,-4,12,1,-19,7,-23,7,-20,4,-8,19,-18,-7,-30,10,4,-23,27,-65,25,-10,-34,7,-4,-15,38,-3,-12,23,0,6,24,-14,-96,-11,46,25,25,38,7,19,0,13,6,12,-22,36,-11,12,-22,-12,42,8,-8,13,-19,12,10,-30,31,-4,-21,22,24,-34,14,-15,19,23,-16,-25,20,18,41,53,7,-24,10),
	(26,-81,0,-19,-31,-8,4,19,-18,19,-68,8,-40,-3,-4,-28,40,-22,-25,27,-7,11,-18,40,25,10,52,-51,15,27,-18,-19,3,-3,13,49,-3,6,15,31,0,9,-2,-13,12,63,15,42,39,15,31,53,-3,7,13,-6,7,-18,7,5,-22,8,1,0,53,6,-14,0,-55,24,-18,-48,-5,18,-1,41,23,-30,-4,41,48,-16,14,-89,-1,61,33,41,19,14,22,4,-13,-1,-2,-19,46,-34,31,-35,-46,29,-24,24,30,8,-17,-22,5,19,-13,-31,11,15,-9,-4,18,-9,34,2,-40,0,6,18,65,23,-55,17),
	(27,-80,-1,-19,-11,-18,-37,3,-12,-30,-57,-22,-32,3,-62,-10,46,-22,-44,-18,-5,-3,-39,49,-17,-6,16,-67,10,18,7,-11,17,-7,-9,23,-25,28,-2,-8,-21,29,-15,0,11,11,42,31,42,37,33,13,-3,0,-28,-19,17,-17,-22,-3,33,-17,-22,-2,41,5,15,-2,-47,-5,3,-35,56,-14,14,52,13,-17,-13,2,28,4,10,-44,25,20,6,35,-7,46,0,15,-5,6,-5,12,44,-14,48,-5,-25,-1,8,40,9,22,-13,-58,4,-27,23,-44,8,13,-39,-32,9,-6,19,2,-28,8,-10,-77,32,-4,-36,25),
	(-4,-23,-7,-10,14,-31,-20,-1,28,-49,-43,-37,-17,30,-27,-50,14,12,-29,-21,34,2,-57,17,-4,31,-35,-4,21,19,24,23,-17,-20,6,21,-9,4,-12,11,-4,13,28,9,2,0,54,-15,-10,38,36,-6,-44,26,2,-29,22,-22,5,-3,47,-2,-45,13,47,1,21,-11,3,-61,44,0,26,38,39,17,-27,-15,-15,-18,5,-18,-20,10,10,-11,-3,32,-46,47,-2,29,0,-5,-7,21,19,-9,10,-26,-38,-37,28,38,33,5,21,-47,20,-19,9,-41,6,11,-9,-7,9,-27,-2,0,-16,2,27,-71,40,1,-24,18),
	(11,-13,9,13,18,-21,-29,6,8,-30,-49,-33,8,21,13,-38,-11,-15,-4,-47,-9,20,-59,25,-22,-5,17,16,27,-17,18,10,8,-3,5,10,-5,18,9,-9,-7,10,27,35,24,-4,14,-6,30,38,0,-7,-23,12,22,-7,23,-22,6,-4,8,3,-44,-11,50,-7,31,-11,6,-69,-1,-22,-10,17,54,-7,-21,-22,7,-6,0,-17,-16,33,-9,-15,-12,-4,-42,12,1,-9,24,-30,-4,44,-38,-12,-16,5,-24,-33,2,-2,22,-2,22,-8,5,-16,-4,-32,19,2,10,-32,6,-43,28,-12,-21,-22,54,-58,7,0,-42,42),
	(-19,16,-4,-2,40,-1,-26,-26,37,-15,-43,-25,14,-3,35,-34,9,-29,-5,-41,-8,21,-14,0,-28,4,-19,3,27,-47,2,43,-19,-7,15,5,-15,1,-7,-5,-21,12,26,11,-12,26,2,42,-6,2,3,-28,5,5,24,12,17,-12,14,5,15,19,-10,-9,69,-2,6,-6,-2,-40,17,-8,-12,8,42,-6,-18,2,29,2,-22,-23,0,20,4,25,1,0,-20,-23,12,11,41,-42,20,1,-29,41,-38,42,-23,-32,-16,-11,-17,-16,-6,-9,24,-24,-2,-44,22,-2,9,-45,0,-20,6,-36,0,-31,50,8,13,-12,-30,25),
	(-13,17,-14,-24,1,-15,-2,-16,26,9,6,-23,24,-1,18,-23,11,-4,-12,-20,0,5,19,-10,-19,-7,4,13,-27,-39,-17,30,-7,22,-34,9,-40,-12,-7,-9,-20,7,38,36,15,-5,-14,-4,17,2,13,-21,20,-2,33,-10,10,-23,13,13,12,-6,5,11,52,12,-14,-7,-12,18,0,-20,-19,33,31,7,2,10,-9,2,12,17,4,5,19,8,-3,12,12,-64,-15,2,29,-47,0,8,-45,30,-17,62,-2,-20,2,20,0,-19,36,-5,17,9,-8,-17,-5,24,-8,-13,7,-12,-12,-14,3,-6,30,34,-3,6,-30,12),
	(-20,-4,1,-1,-43,-25,-4,-5,-12,13,18,-9,-8,19,0,-28,5,-7,-30,6,-3,1,15,-20,9,-15,0,31,-9,-16,-7,38,14,7,-27,26,-27,-13,-30,27,12,4,16,28,18,-8,3,23,-9,6,-23,8,-5,18,25,-6,17,21,24,15,16,10,-12,9,0,19,-6,-16,-11,11,-9,-22,-11,46,5,8,11,3,15,-21,-18,13,-7,6,3,52,30,-10,3,-46,1,-18,25,-14,21,10,-58,-3,23,57,-31,1,-23,15,14,-10,1,-3,9,16,19,-21,-5,11,20,-6,-3,25,2,8,-14,-32,-5,12,24,26,-2,27),
	(-45,7,-10,13,-54,-13,9,-2,0,-5,10,-7,16,45,-2,-33,-30,-10,-29,-19,3,10,-17,-6,7,6,-11,13,-16,-48,1,30,39,-3,-56,22,-13,17,1,-14,2,14,6,51,28,-38,21,7,-10,-23,-5,38,-3,16,-3,3,-20,17,9,0,0,-26,16,33,-26,-2,-16,13,4,11,-9,-12,-27,3,19,-23,16,10,18,14,-21,23,4,-21,16,28,32,-34,7,-19,-10,5,2,6,17,-5,-38,6,-17,46,16,16,-5,20,-14,10,14,23,12,7,15,-3,8,0,35,4,0,-13,-1,8,-49,-21,-17,2,9,-12,-42,-9),
	(-64,10,1,18,-29,2,0,-7,-9,-11,-19,0,-16,1,17,-3,-17,-11,-22,-11,-15,28,-14,13,-12,-7,-9,36,-8,-41,-13,13,4,-10,-3,0,-36,-8,16,-25,12,51,-14,6,23,-15,35,-9,13,-7,0,10,-12,13,-9,20,-18,21,1,-17,15,8,24,-4,-37,29,-23,-16,-30,0,17,-19,-37,-29,15,-30,9,18,14,-11,15,26,-15,4,15,16,53,-45,23,-4,-27,3,-6,6,14,-9,-22,3,-5,52,18,4,-23,5,-11,26,6,13,33,-7,21,35,-4,24,11,20,13,-6,28,-12,-49,-2,-41,20,4,-11,-22,-16),
	(-44,-6,-1,32,5,1,41,-28,-5,-31,-21,-29,-35,-18,37,-8,2,-13,-3,-37,16,55,6,38,-13,16,22,-17,-13,-29,-22,44,5,-31,-3,-17,-44,-47,-11,-31,-15,9,13,2,0,-21,14,41,-6,19,0,-4,4,-12,-42,31,-26,10,-3,-11,12,-7,11,7,-54,-7,-31,19,-31,-24,31,-16,-31,-34,-14,-10,1,15,13,15,8,19,-21,22,5,-5,43,-50,1,-7,7,-16,9,16,19,-15,12,-11,-51,1,14,32,9,2,18,27,-8,43,19,-14,-3,28,-8,-23,18,36,-9,-28,6,-24,-76,16,-15,11,20,3,-40,-1),
	(-92,0,-8,-2,-17,-11,25,-39,-12,25,-15,-20,-37,-56,10,-4,8,0,-23,-16,21,53,23,20,0,5,4,2,4,-19,-39,52,-9,-40,1,-44,-63,-31,-1,-38,-3,10,0,-47,-38,-28,18,-1,-1,34,20,-27,22,19,-1,-14,-45,-12,29,9,19,-4,-16,7,-42,10,-6,-2,-16,-2,-15,-27,-29,-55,18,5,-1,1,28,6,8,-31,2,-23,-7,-11,34,-49,-14,6,-7,2,33,30,1,3,-14,7,-51,-12,24,23,33,-12,11,15,12,36,24,16,8,29,10,-27,25,38,2,-33,4,-37,-62,12,-35,25,20,-19,-35,-2),
	(-93,47,-19,-4,0,11,38,12,-4,17,-49,-3,-30,-57,-1,-14,-8,-14,8,-12,43,20,6,43,12,-13,-33,0,10,-1,-52,33,-9,-23,-7,-24,-79,-44,26,-72,9,1,-20,-33,-29,-4,-10,2,-12,21,-4,-33,34,13,-23,13,-30,3,12,-2,20,-34,-49,1,-55,33,0,18,18,-25,14,-56,-26,-40,23,-7,0,-18,-6,6,27,4,-9,-19,-28,-35,-4,-43,-14,41,-12,31,57,27,16,-16,-7,22,-68,-53,19,47,37,-17,14,40,25,28,9,-26,27,42,15,-61,1,18,34,-30,36,-16,-83,-4,-50,-38,-9,23,-55,10),
	(-75,28,-33,-23,-17,0,26,24,10,32,23,31,-10,-24,-19,3,1,27,-3,12,-18,-9,15,5,5,14,33,-8,38,3,-25,16,-12,-22,12,-14,-65,-33,-2,-90,-17,0,-40,-35,-20,-7,40,27,-45,-37,44,-20,24,-61,-45,-30,-46,-5,-21,21,-24,7,-31,2,-47,-1,-7,37,14,-16,30,-31,7,-23,-26,11,20,-33,-32,52,4,-37,-4,-16,-10,-41,-50,-40,-49,-33,-51,16,25,7,-50,-57,-1,35,-86,-44,27,47,-19,13,21,48,-34,-16,2,-32,-8,17,20,-52,-23,41,60,-37,37,-54,-95,7,-13,-4,8,8,14,-20),
	(-59,-26,10,-6,-2,-21,-11,15,28,-24,31,30,-10,9,-26,3,-16,28,27,-2,18,-26,-30,-46,-14,3,7,-26,10,-4,-3,21,-18,-26,54,-11,-17,14,8,-33,-31,4,-15,-36,-22,-2,20,30,15,-19,21,14,-21,-23,15,9,-10,-16,-35,-17,-19,-11,6,-68,-22,-18,54,14,27,0,-4,14,14,-4,-36,4,22,-27,-20,19,-30,7,-17,8,1,-16,-12,-48,-66,-18,-57,-32,44,-18,-32,-34,28,20,-24,-53,23,-8,-42,-11,39,28,-13,-23,-7,-61,-21,-17,-21,7,7,-33,8,9,-8,-13,-37,6,13,1,-11,-29,10,-6),
	(-28,-23,41,-25,-19,-48,-37,-25,-1,-40,37,18,-6,1,-26,9,-38,19,-15,5,65,0,-22,1,28,8,0,-18,1,12,25,-25,24,9,44,-24,-8,39,-33,20,-3,27,10,-39,2,-27,11,19,33,-29,-11,14,-11,41,39,30,-8,-1,-30,3,28,15,-17,-43,-61,11,59,-33,6,27,-10,-17,55,-24,-15,-13,20,-4,-55,-7,-34,18,-35,-10,12,-26,22,-11,-40,8,-30,-30,49,-42,-7,-25,-10,28,6,-12,1,-5,-44,1,26,-6,-11,-30,-18,-23,-3,-4,-39,-24,12,-35,-40,6,18,-14,-8,-5,0,-30,-4,-40,-14,-2),
	(-47,0,-1,5,-28,-22,37,-4,15,-12,-4,-9,6,26,3,2,-7,2,0,-2,32,-9,-22,-12,-4,-25,-48,-4,13,-5,4,3,-14,-15,31,-5,6,12,-34,7,-20,0,44,-20,-12,16,20,-8,13,20,1,-30,3,37,2,13,-5,-1,18,10,-5,3,-4,-16,1,15,-22,-46,-15,-16,-21,-6,28,-23,-1,-4,-16,-26,23,-24,-39,-13,-10,48,-11,26,7,-22,-22,42,-2,-20,19,-15,26,-42,6,28,-16,33,-32,-15,-27,-17,28,-6,-17,24,-9,17,11,-10,-45,-12,17,10,-38,12,-43,-14,-21,-20,25,-10,19,-4,3,1),
	(1,-11,-15,12,-6,2,9,-4,0,12,25,-2,-13,19,-21,12,-10,-12,9,2,13,15,3,18,15,-2,-12,-7,2,26,0,-4,-7,-6,-12,-7,-8,6,-1,-9,-7,8,4,4,-23,1,-12,11,5,-2,-17,-19,2,4,16,-8,9,-4,-7,-10,-23,8,-20,15,29,9,-13,8,-23,-3,23,12,-7,-4,10,2,-3,6,-3,-23,-10,-17,-2,5,3,15,0,14,11,26,14,-16,2,21,-8,-14,-10,-20,5,-4,15,15,-23,9,-10,17,8,-16,-17,14,-21,-3,-10,-20,-20,-5,-4,-13,8,-7,-7,-15,-8,-20,20,16,2,-6),
	(12,-15,-7,-23,-6,-16,-15,-19,-2,3,37,0,12,-5,18,23,-6,-8,-10,-6,34,22,29,0,17,-23,-9,-17,16,24,7,20,0,-20,20,-13,21,-18,-20,6,30,-2,20,-21,-32,17,-8,18,6,-9,1,-22,39,4,10,23,-9,23,7,-3,-10,-8,-7,-23,-10,16,0,-24,25,33,-38,-4,25,10,-21,-17,1,-10,3,5,9,-18,-26,10,-10,35,2,-31,5,21,19,-19,17,7,16,-27,0,-7,8,40,19,5,-4,-11,8,19,-15,3,8,17,-7,-7,-9,28,-5,-28,-30,0,-15,13,23,21,-26,33,0,4,12,-33),
	(8,-17,13,-35,3,-36,4,-29,8,31,45,9,34,8,12,2,4,19,32,2,20,32,-8,-6,23,-38,-20,-30,12,-2,-44,9,-43,-22,35,-14,18,-21,-5,4,23,49,42,-22,-27,13,7,-21,33,12,19,-35,22,-15,30,10,-14,-2,30,-7,9,-2,-9,-34,-41,23,-15,-3,23,33,-48,-9,11,44,-9,-23,-44,-8,33,-1,-5,-34,8,32,-10,35,5,-32,-23,17,-5,-31,7,4,19,-33,-27,-23,6,53,-16,-7,-15,-10,7,-28,-13,-2,-22,7,14,-1,-14,22,6,-17,-38,3,-20,16,-1,5,14,38,3,-18,8,-42),
	(7,8,-1,33,21,-1,-9,28,13,8,-39,27,11,25,6,-2,-40,30,-31,-25,-13,20,0,-34,8,-2,-20,15,-2,21,7,33,-7,-24,-1,-26,-28,16,-18,2,-3,11,40,-3,-9,24,5,-9,13,-6,-1,8,25,17,18,14,-7,-38,29,9,2,-35,-11,-34,7,-12,25,-51,-72,2,-3,-7,2,32,-24,-32,-23,2,-15,-32,-36,3,-18,6,23,-3,6,-30,-32,26,-33,-23,34,-3,33,-30,-18,-8,10,26,-30,-28,-8,1,5,8,11,20,-23,3,20,31,-17,-1,21,-3,0,-5,-34,10,-24,27,32,46,-17,-1,-19,7),
	(-1,28,26,4,-14,-32,6,19,-51,-8,2,8,-44,12,4,-37,-17,-16,-44,-37,-11,37,23,-31,40,1,-8,-27,-11,1,-10,23,-6,-4,-17,-6,-11,-10,-18,-26,25,34,30,-20,-17,-14,-29,-35,16,0,-41,-32,-15,-4,-33,26,-15,-45,25,-14,17,-69,-49,2,-5,14,18,-31,-79,-45,3,-20,3,25,-11,-32,-22,0,8,-29,-15,27,-6,-8,-6,-34,12,-23,-29,-8,-16,21,20,-17,40,4,-22,-7,-16,46,9,-15,31,10,-20,-7,46,0,30,-4,32,41,-2,-21,-25,17,-6,-9,-44,-36,-37,-13,39,-6,-16,-29,-43,27),
	(2,28,31,-1,21,-6,3,41,-55,8,12,26,-32,-30,8,-58,3,-16,-55,-50,3,-4,8,-14,15,-3,17,-19,-5,24,2,10,6,-39,-9,-29,-2,-36,-6,8,-4,-4,4,-16,-9,-3,2,0,22,18,-39,-1,16,13,-29,17,-42,-22,37,-2,20,-33,-49,-4,-89,35,2,-1,-103,-12,13,-29,31,-26,20,-12,13,-11,-10,3,3,0,-14,-21,-21,-13,64,-11,-47,9,-37,18,20,-14,29,-11,15,3,-13,4,27,20,-18,10,-37,17,2,1,-27,-12,11,27,13,-13,4,0,-7,-9,-44,-27,-46,-19,-7,24,-25,-26,-45,4),
	(36,25,39,9,24,16,30,8,-61,61,-19,47,-24,2,16,-42,14,4,-10,-34,-15,25,44,-7,20,3,12,0,-15,-10,-30,8,-18,-45,-4,16,-9,-23,-26,-18,7,-28,-5,-33,20,8,-26,10,11,14,-11,5,-4,4,-37,2,-37,-23,18,11,10,-32,-42,15,-28,7,-6,1,-61,-4,6,-5,32,-12,9,10,-2,-8,9,-1,4,18,20,-30,0,-30,38,-37,-2,24,-17,0,-18,29,-4,-15,8,-14,-22,-6,-3,31,-2,10,-19,27,4,-5,-18,-2,2,20,-2,-4,-8,-3,3,8,-9,-15,-19,-6,-23,51,-3,1,-19,14),
	(14,43,60,-1,6,24,2,9,-61,62,-38,46,-40,24,0,-18,-5,13,-13,-27,11,25,12,-43,10,3,29,-8,-44,-17,15,-1,-1,-13,-10,7,12,-12,8,-22,11,-18,-55,-15,7,9,-57,9,25,2,-32,-1,21,3,-15,6,-38,-1,31,-5,-12,-11,-10,32,-8,36,-10,8,-105,31,9,-6,34,0,7,30,19,-10,-9,-5,23,21,12,-8,-15,21,45,5,10,-26,-3,17,17,9,12,-26,45,-20,-54,-15,21,30,-1,16,-38,-9,12,17,-11,15,4,1,5,-34,-37,-5,-40,-28,9,-3,-11,2,-35,23,-10,31,-31,32),
	(0,32,53,16,-2,26,31,-23,-12,58,-21,24,-9,9,11,-44,-21,-22,-4,-17,18,26,15,-43,-7,-7,7,-16,-4,0,-1,7,-22,0,-20,19,-14,0,18,-11,-8,-9,-42,2,-5,-9,-42,-3,-1,-14,7,17,6,-14,-13,2,12,3,4,-1,-8,18,-27,21,-6,17,-13,4,-90,19,-14,-21,-5,4,-20,17,-8,5,4,-1,16,-6,12,-27,-5,7,38,10,21,-10,8,20,-4,15,19,-10,1,-17,-51,-19,9,35,12,16,-31,-1,16,0,-6,12,5,-35,27,-2,-1,18,-3,-11,20,-37,-32,-19,-1,29,-3,-15,-35,2),
	(1,2,45,4,14,27,-10,-32,-23,62,-32,22,-28,-14,16,0,8,8,0,-30,-5,45,12,-12,-1,-28,39,-10,-17,10,-12,-32,-17,-21,-3,19,0,-17,0,9,-13,18,-51,0,-1,21,-24,3,32,-8,16,0,4,-7,2,-18,-4,-17,17,-1,-19,10,-2,5,0,34,1,2,-96,41,-15,-8,-1,0,-13,19,7,1,-7,-11,29,-6,12,-59,15,7,9,35,32,36,0,5,20,9,27,-2,3,-8,-10,-8,31,43,24,0,-22,13,2,-20,-17,-3,-3,-33,26,-2,4,0,-14,-6,3,-20,-48,-16,-6,46,-1,32,-2,26),
	(4,-28,20,-17,-12,10,9,-18,-22,47,-87,29,-36,-29,15,-13,33,-35,-35,5,-19,22,-26,8,19,-36,20,-18,7,14,-15,-33,5,5,-11,-12,20,-11,17,0,5,8,-36,5,36,46,-49,-8,18,-5,29,22,19,-31,0,6,34,1,14,-4,3,36,26,0,13,11,2,21,-48,16,-22,-28,4,-12,0,13,6,-25,5,-9,16,35,10,-70,-32,17,25,14,31,20,39,-21,27,-13,-2,10,16,0,33,-17,12,49,8,-6,-29,-10,13,13,11,22,-13,-23,18,-17,-21,14,13,-22,6,-18,-7,-14,-23,39,48,41,-23,19),
	(22,-71,9,-26,-15,-15,-17,0,-14,39,-103,33,-42,-28,28,-8,29,-20,-24,8,-33,0,-28,0,1,-16,31,-47,-11,21,3,-25,12,1,-1,12,16,-9,37,-2,-11,12,-33,7,28,23,-27,16,13,-15,44,50,11,-16,-25,-10,-1,-9,-6,-20,-25,23,41,-4,22,31,14,16,-36,26,-16,-48,7,7,5,35,0,-35,14,4,11,36,-18,-39,-17,34,30,33,16,23,20,18,3,9,8,-10,29,33,14,-14,-8,25,-20,-13,2,21,-16,-21,10,47,3,-31,13,36,10,-4,-14,-22,13,-36,-44,-9,-9,-3,38,17,-22,7),
	(36,-88,-9,-8,-14,16,-15,21,-1,-26,-90,35,-63,-11,-30,22,25,-7,-60,6,-30,14,-35,17,36,23,39,-37,20,18,-10,-11,21,-1,-28,29,-14,29,31,-8,-21,-5,-23,-12,22,-14,17,50,23,8,30,24,-12,-30,-1,-23,5,-38,0,-8,-13,21,25,11,32,7,-2,-2,-25,-2,23,-43,13,-16,18,39,18,1,-20,20,23,26,-22,-49,-13,24,39,8,4,32,19,13,-16,-1,-9,11,10,1,38,-28,-7,23,13,12,-7,32,-1,-30,11,19,-6,-35,29,17,1,-1,-10,-8,42,6,-16,33,-27,-56,37,21,-20,-1),
	(37,-59,-17,16,-8,12,-14,0,30,-56,-28,2,-52,15,-20,15,13,17,-36,-5,-21,9,-55,15,-12,46,18,-7,25,30,7,-6,27,-4,-23,21,12,15,38,-4,-36,0,25,-4,52,-7,33,37,21,13,-3,18,-28,9,-3,-9,15,-24,-20,9,23,32,-11,22,40,7,-14,29,14,-54,36,-8,13,-5,43,21,-4,22,-25,-2,21,36,-20,5,25,4,7,28,-19,35,-18,7,-11,-21,-8,45,28,2,51,-7,-13,7,22,15,21,25,5,-19,34,-30,4,-46,24,26,6,-18,23,-22,41,-6,-11,23,-19,-106,9,-18,-12,26),
	(47,-26,-14,-8,-15,13,-19,-7,19,-21,0,-9,7,56,-5,-26,0,0,-10,-22,6,13,-47,14,-9,12,-26,1,39,6,22,18,18,-2,19,52,7,8,0,1,-12,27,45,8,12,-19,67,0,-2,14,5,5,-13,0,28,-4,25,-22,-6,0,14,22,-3,2,74,-1,24,4,18,-34,26,-5,-6,24,53,12,5,24,-28,-16,-6,4,-37,49,-6,-19,-1,18,-21,31,-27,14,4,6,-25,36,8,21,12,-5,-2,-15,26,38,0,-10,12,-25,9,-19,28,-10,36,4,-16,-8,0,-20,29,-6,-8,-5,26,-79,10,-24,-24,15),
	(14,0,16,-13,6,33,8,16,26,-23,-36,-8,-3,27,3,-28,-32,21,-17,-45,-21,-5,-57,19,-10,9,-7,7,21,-35,8,9,-33,19,5,49,2,31,9,-13,-8,37,51,0,25,-21,17,31,-11,11,20,14,-13,6,22,23,14,1,-7,-19,9,14,-16,21,57,0,-10,24,-10,-32,36,-2,-42,-4,39,0,-4,-8,11,-20,19,5,-19,43,2,-3,-13,-11,2,-20,10,-5,0,0,4,20,-28,43,0,16,-27,-8,-13,20,5,3,13,10,3,-21,13,-46,13,35,3,4,4,-49,16,-5,-19,-7,29,-30,14,-11,-10,23),
	(36,-15,7,-4,38,13,8,12,34,-18,-42,-36,-14,17,3,-19,9,-8,6,-19,-17,1,-7,10,-16,16,-2,11,-11,-24,9,35,-24,9,13,43,-26,4,20,11,-8,-19,29,31,21,11,17,0,14,-3,31,-38,12,2,12,0,28,-22,5,14,-4,9,-7,3,24,-11,13,-12,-16,-13,0,-8,-39,7,21,12,19,-2,35,14,10,0,-1,8,-3,41,-29,-6,27,-1,2,7,-30,-35,-8,24,-31,41,-5,48,-3,-24,-15,2,-3,7,18,38,27,3,11,-29,2,15,1,-17,4,-10,-3,8,-5,-21,56,6,-7,3,-34,30),
	(8,14,1,-14,8,-8,-1,-26,10,-16,0,0,-1,10,11,-38,-6,-13,-17,-5,-1,13,-16,0,-15,9,-1,1,-2,-16,-3,21,12,-8,-25,25,-12,15,-8,24,15,-30,10,31,25,12,-5,22,1,13,8,-29,-1,7,27,10,15,-14,23,-13,-12,-16,-9,4,48,7,0,-11,-6,-14,12,-13,-14,9,31,-7,8,8,12,0,-13,-4,12,13,-6,37,4,-5,13,-28,13,0,-31,-46,1,18,-18,26,1,20,-10,-3,-11,8,-12,4,17,-3,38,0,24,-23,6,7,26,-33,-3,11,4,11,-13,0,27,21,7,4,-45,5),
	(-15,4,-18,10,-34,0,15,-18,7,-19,3,4,-7,32,0,-10,6,-14,-42,0,-25,21,-3,0,-32,-24,10,4,-19,-38,7,26,5,23,-20,14,5,-9,1,4,-23,6,28,44,29,12,17,2,4,-2,15,15,5,-18,16,32,7,26,31,-6,0,-12,16,16,-18,0,-40,-10,-4,-9,-4,-12,-9,34,-1,-3,16,7,10,7,-6,26,-6,4,-9,56,28,19,31,-30,0,-15,-32,-18,5,-1,-8,22,30,42,-13,-2,5,10,-19,6,33,28,14,14,15,-23,11,6,24,-18,13,17,-5,-6,9,-7,-10,-1,16,-5,-27,25),
	(-4,-3,-31,15,-29,-13,18,-12,-15,-12,-10,-22,8,6,-5,-13,-4,0,-17,-25,-41,3,-50,7,1,20,18,1,-6,-27,-6,13,34,41,-17,-37,-20,-25,-14,-4,-6,39,-5,39,18,-9,14,33,-3,2,-5,19,-15,-5,-14,15,9,-6,22,9,-8,-13,-9,11,-45,12,-43,-13,-13,-19,-3,-38,-27,-3,-5,-6,16,23,-11,-7,-18,20,-11,7,9,33,18,9,24,1,-23,-26,3,-17,21,9,-25,42,5,14,-1,19,11,-10,-36,9,24,50,32,39,20,24,23,20,16,27,0,19,19,5,1,0,-36,-18,29,2,-36,14),
	(-27,-3,9,-2,0,-3,36,-13,-1,-8,10,-22,-5,-7,35,-29,8,5,-21,-32,-11,14,-47,0,-2,-10,8,-1,-2,-45,5,7,-3,13,-15,-33,-16,6,6,6,6,36,0,-11,24,6,29,3,24,0,-15,21,-7,6,-13,37,-5,-21,25,-12,-7,1,19,8,-60,0,-18,-9,-8,-28,-9,-29,-38,-45,21,-4,-1,35,26,8,0,21,-9,13,-9,28,33,7,16,21,-22,-22,-7,10,-3,2,-21,17,7,44,-13,23,-10,-3,-26,10,1,36,19,7,28,30,-1,-12,7,6,-16,8,20,1,4,0,-49,1,10,-18,-46,-8),
	(-64,35,10,0,19,-11,24,-30,2,0,5,1,-16,-39,43,6,24,-32,3,-28,6,18,-23,33,2,-12,28,5,-17,-52,-26,17,-1,-31,13,-46,-5,2,-24,-27,-6,36,6,-14,1,0,1,4,3,6,15,-21,-11,-4,-23,-7,-25,0,4,14,-16,-2,13,32,-64,19,-53,-24,-15,-11,20,-20,-37,-11,14,-14,1,10,32,-7,13,10,0,27,-10,9,52,10,-11,20,-6,-1,-9,22,0,-11,14,10,-6,23,29,39,11,-37,-2,20,1,46,13,18,22,31,-2,-23,22,16,10,-24,-11,2,-31,-11,9,3,16,7,-37,-1),
	(-73,18,0,-2,26,0,20,-4,0,-4,-16,7,-40,-66,15,-12,11,-34,-33,-8,7,38,12,40,21,-20,-2,-8,-15,-53,-39,-6,-9,-13,-4,-14,-21,-28,-17,-30,-5,-19,37,-9,2,-3,-7,1,-22,-1,24,3,14,15,-28,18,-44,3,7,7,14,11,-30,15,-68,24,-49,-11,-39,-20,9,-30,-58,-38,-6,-3,6,7,4,21,12,-6,17,12,-6,-26,30,-21,4,16,-12,-11,0,15,19,-27,16,26,-44,-22,9,31,18,-29,17,14,11,20,17,-8,-14,34,15,-42,-20,12,-8,-35,-18,-14,-40,34,-6,-7,-10,7,-39,-24),
	(-67,39,-23,-31,2,19,35,3,-9,0,-22,-6,-7,-44,0,-2,7,-13,-44,-17,3,20,0,34,-2,20,-27,-18,35,4,-24,22,3,-7,10,-5,-39,-36,-30,-42,-9,-5,30,-17,-9,8,33,18,-32,0,29,-12,28,12,-19,-28,-38,-36,-4,-5,-21,-36,-43,-7,-49,7,-50,48,-13,-17,29,-59,-27,-29,3,6,-24,-47,-6,37,5,11,26,4,-15,-18,30,6,7,34,-18,-11,26,33,-31,-66,7,12,-81,-61,48,37,27,-40,32,36,-19,17,-12,-16,-39,15,29,-28,-46,43,34,-40,-23,-24,-54,2,-17,-11,42,20,-1,-30),
	(-80,0,-2,-16,-32,15,18,-14,25,42,4,30,-38,-33,-21,8,31,-6,-16,1,11,-20,15,10,2,30,-20,-20,0,-9,-21,12,3,-18,-7,-23,-40,0,-22,-64,16,-25,4,-10,-21,-11,24,24,-39,-53,22,-13,24,-2,4,6,-42,-32,0,13,-30,-16,-22,-30,-17,-11,-60,6,70,3,7,-50,-63,19,-7,42,-9,-6,-4,25,-35,-48,9,-18,-22,-24,7,-29,-29,-8,-14,-37,40,31,-46,-66,53,19,-81,-35,11,-9,-52,-39,40,31,-33,15,-18,-16,-48,-3,-7,-24,-25,28,43,-13,1,-4,-74,17,36,-8,31,5,7,-37),
	(-72,11,17,-6,-4,0,8,38,18,31,-12,10,-34,21,-33,24,15,12,-19,29,13,-23,-1,-15,-24,-12,3,-9,16,-1,-1,-23,-24,-26,28,-32,11,23,-31,-42,-44,-17,10,-26,-31,-23,10,10,-7,-51,-1,7,-14,-8,15,36,-37,-9,-37,20,-38,4,16,-39,-25,-36,-9,-8,43,-19,-17,-6,-16,4,-33,0,5,-38,9,31,-27,-21,32,13,-19,-1,1,-33,-58,-10,-52,-15,-14,3,-2,-21,49,23,-40,-18,28,-19,-49,-12,22,11,6,-9,-2,-14,-12,-27,-37,-17,17,-11,-23,0,-13,-46,-40,39,15,-21,32,-8,11,-8),
	(-30,-52,-6,12,-6,26,22,-7,10,-7,46,-17,9,-12,-9,3,2,-3,-18,20,3,-28,-23,-30,-33,32,15,-11,34,-6,31,-28,-4,-4,28,-12,0,33,-30,1,-20,-17,11,-4,-3,-32,3,1,-1,-16,1,23,-10,8,49,69,-49,-15,-39,-15,-17,35,21,-15,-54,-9,21,-28,51,17,2,2,2,-12,-50,2,71,-18,-20,9,-45,14,14,-11,13,-4,25,-11,-57,-9,-38,-34,-18,-31,-15,-31,-1,41,-15,27,25,-10,-43,-17,12,22,-4,-37,-15,-19,-8,20,-37,-25,28,13,-2,-3,-8,-25,11,10,41,15,16,-50,9,-6),
	(14,-23,-8,3,0,33,0,-16,38,-13,9,-12,5,-21,-3,22,-8,-3,28,15,34,-17,-7,-7,-31,43,3,7,9,-25,43,-13,-10,-3,39,-19,-8,43,-12,-39,6,0,30,28,9,-29,-5,24,-24,-4,27,6,0,12,5,22,-10,2,-21,0,-32,4,8,6,-16,0,-4,-18,0,-4,38,-8,-39,8,-18,4,10,5,-21,26,-28,13,22,-35,-14,-11,-5,31,-31,-23,-29,-8,-16,26,-23,-1,6,26,-2,-8,30,-20,9,23,0,29,9,0,2,-11,9,21,11,0,14,37,29,16,-12,-6,-9,42,17,-17,15,1,12,2),
	(-15,8,-8,-15,-17,-18,15,0,-5,14,-5,14,-13,5,-10,-6,-2,24,-5,24,13,17,-19,-10,-15,0,-2,4,6,-8,18,-27,-14,6,-8,-1,2,1,3,-3,-6,7,-25,-1,-6,6,-13,9,16,12,-5,18,20,-18,-5,-18,19,11,-10,13,-13,3,0,9,5,12,-14,10,16,-2,-21,22,-5,8,-3,-21,5,-12,5,-8,-14,1,7,-10,14,13,2,-13,8,8,13,14,12,15,0,-21,-12,-15,30,-20,-2,17,-12,0,22,-13,0,-8,-9,14,-7,-1,15,10,3,7,-6,20,-3,23,8,23,2,3,7,7,13,-27),
	(-12,-6,6,-4,-9,-21,6,-2,-6,-1,-5,23,-3,15,0,0,12,-27,8,8,10,15,-5,-22,15,-24,9,-31,9,-1,-3,-7,-4,-10,4,20,15,14,0,31,23,-13,23,14,12,8,14,-5,12,25,-2,0,29,12,1,-13,6,14,20,-1,29,-34,5,2,-6,-5,11,29,21,4,-1,18,30,21,27,-13,-15,-7,-7,16,-21,-5,-10,1,-12,4,2,-10,9,5,-10,13,13,2,-19,22,0,6,28,29,-4,-27,-7,-21,1,-21,16,12,20,-27,17,-25,0,21,20,-38,-13,29,21,-2,-7,-11,0,23,16,-23,-26,16),
	(-2,-43,-13,-3,-13,-35,-25,-56,24,23,24,-13,29,38,21,10,-29,26,20,29,30,67,-1,5,34,-10,-11,-34,1,-10,-18,54,-30,10,17,-13,2,-6,-11,34,39,34,37,19,-23,17,-6,15,13,33,3,-22,43,8,8,4,-21,31,13,-10,23,-10,-11,-7,27,25,-19,-33,1,6,-42,0,11,12,-10,-16,-21,-16,19,11,2,-24,-20,33,-47,11,8,-8,-29,14,28,-16,17,8,-15,-5,-18,-26,9,58,-6,-23,-11,-49,9,-27,-18,20,-9,21,-13,-43,-32,21,-2,-34,-40,3,0,33,17,-14,-2,60,30,-20,9,-11),
	(-15,-31,0,15,-2,18,4,4,-25,33,-30,-17,4,36,10,-8,10,9,-8,11,12,11,-23,-26,6,14,22,4,10,19,31,35,-13,-32,9,-24,6,-17,-34,-4,-8,-5,18,-3,-4,22,-30,7,-6,6,-20,-22,-16,12,29,7,-28,9,-18,0,5,11,5,6,-14,-15,9,-33,-58,8,19,-15,31,30,-7,-22,9,-19,-23,-27,-15,-15,22,33,-1,16,26,17,-14,33,-1,-19,-6,-29,20,-29,15,-7,18,3,-3,-41,-34,-5,-3,-24,9,-27,-25,-27,19,21,-18,0,17,-10,-17,17,-9,-6,-10,-5,14,13,36,-19,-1,4),
	(0,33,11,-1,39,4,-5,28,-28,0,-15,-13,-71,2,20,-13,-6,-16,-1,-25,-23,-5,20,-34,-7,-19,22,-18,0,23,-2,-17,-14,2,-41,-32,-2,-10,2,-1,19,20,8,-44,-6,13,-28,-15,11,-1,-55,14,-3,2,5,24,-21,-28,17,-16,-9,7,11,-2,-12,34,-21,-55,-72,-4,-34,-20,-1,15,-28,-34,-10,-13,-8,-18,-3,19,-5,31,-7,-16,19,9,-41,1,-1,3,0,8,23,8,-12,-15,-4,9,23,-28,-1,-21,-47,-22,0,-4,7,-14,26,47,-7,9,-31,14,-21,-9,-29,-19,-27,10,14,-12,-21,3,-11,1),
	(5,20,18,-11,19,5,-6,10,-63,31,-70,8,-54,-29,8,-40,11,-22,-13,2,1,14,32,-8,23,-34,13,-21,-2,-20,-35,-13,-21,-49,-25,-9,7,-48,-19,2,-12,-16,-10,-57,20,-5,0,29,19,5,16,25,-5,-18,-46,5,-40,13,36,12,4,42,-23,-9,-54,26,-6,-12,-100,0,-20,-48,51,-23,-14,-11,0,-3,16,26,-4,4,-6,-35,-9,-9,25,-14,-47,14,17,-29,-3,38,-11,-13,5,-15,-38,-2,10,36,-8,-11,-33,14,13,-9,-4,-6,5,1,5,10,-26,34,-15,-24,-28,-40,-36,-3,-2,30,-13,-6,-48,-2),
	(46,46,36,0,13,20,11,23,-47,59,-52,25,-16,21,26,0,10,12,-20,-28,1,6,6,-42,-3,10,13,0,-34,-2,7,7,-19,-33,-2,-21,-20,-11,-26,0,-14,13,-30,-57,5,18,-26,43,-18,-20,24,31,14,-38,-60,-19,-35,-21,10,-3,-17,71,-28,18,-70,-4,31,15,-81,31,23,-32,29,-4,-4,13,-7,9,-16,13,5,0,25,-56,3,-3,43,-7,-15,-13,-11,-23,0,-1,18,-31,17,7,-22,-13,41,13,-28,13,-46,22,22,7,-4,11,15,-6,0,-12,-14,-4,-9,-24,-23,-21,-51,-4,-28,17,4,-8,-23,8),
	(7,45,53,-14,7,6,13,7,-52,44,-80,32,-8,14,2,3,-6,10,-21,-12,-13,14,10,-31,27,-11,21,-2,-12,3,-10,-22,-18,-17,-20,-3,-4,-5,-29,2,-5,0,-48,-43,12,-7,-36,16,-10,-23,0,27,20,-37,-14,0,-19,8,27,0,0,42,8,19,-17,29,19,19,-66,9,10,-20,4,-15,-25,37,3,-11,11,-1,26,-6,48,-33,4,22,30,10,-13,-22,-9,11,6,32,6,-25,-8,-5,-61,7,39,21,-15,17,-47,5,16,13,23,28,7,14,-9,-35,-18,-7,-18,-13,-16,-26,-11,0,-21,-6,14,16,-26,-2),
	(14,32,48,4,27,13,29,3,-38,62,-97,29,-18,22,15,-3,6,-7,-25,-6,-11,54,11,-21,-1,2,17,-15,1,29,-3,-31,-25,0,-3,-13,-14,0,23,9,-32,-1,-44,-17,-1,4,-42,11,-3,-4,25,18,21,-26,-13,2,-14,6,22,17,3,14,20,21,-15,25,15,5,-41,-3,6,-17,-7,-5,10,20,0,-14,23,21,26,-5,35,-21,12,20,23,2,13,33,26,1,19,10,0,8,-17,-6,-42,-2,17,45,10,0,-16,12,25,-28,27,23,-5,-20,15,-20,5,-1,-24,-42,7,2,-18,-22,-18,24,14,-7,-17,14),
	(17,-13,39,-19,2,-4,21,-27,-27,16,-122,21,-47,27,13,-14,45,-26,-37,18,-14,52,9,-6,13,3,21,-5,-3,39,-4,3,-36,11,-12,0,-10,-37,40,-20,4,-22,-42,-21,-10,17,-30,13,25,9,18,10,15,-29,-15,-11,34,4,12,17,-21,39,35,10,12,15,1,30,9,14,-13,-25,16,-15,-14,-1,3,-1,4,9,39,-16,25,-29,5,22,37,30,22,24,41,-17,36,25,11,-17,-27,0,24,3,44,22,10,-19,-9,-6,-4,-4,24,15,-5,-19,0,-32,22,30,-13,-28,15,15,-50,-18,3,8,17,6,-31,2),
	(-11,-45,32,2,15,-10,22,-43,-33,25,-89,25,-53,-13,14,24,41,-7,-45,10,-4,19,-29,-27,22,-19,9,-32,16,9,8,-22,1,34,-4,-22,10,-17,29,-2,11,-19,6,9,6,34,-28,18,24,5,56,6,32,-23,-4,-17,18,9,-3,5,-7,29,21,5,6,15,4,29,15,17,-22,-43,-19,-12,0,19,17,-16,0,-12,-4,-13,10,-47,-34,25,5,17,33,14,14,-10,27,12,3,-26,-42,-1,14,-13,53,10,-12,0,4,25,2,-11,29,22,-12,-59,10,6,-7,1,-2,-5,27,7,-31,3,21,2,49,18,-5,0),
	(-18,-67,8,9,-2,27,10,-25,-23,-25,-94,8,-55,-13,9,12,50,-2,-51,4,2,-12,-23,14,13,-14,1,-11,-10,35,6,-18,-4,28,3,1,2,-7,22,-16,-36,-9,-8,-5,22,-3,12,30,16,26,27,18,6,-9,-4,-1,8,-28,27,-1,-4,15,49,29,24,9,-16,29,18,20,-6,-25,-6,-12,-29,36,25,-10,3,7,-5,28,-6,14,4,-14,28,-25,12,18,0,-11,13,-2,-3,-24,-25,33,37,-3,15,28,-8,7,2,6,21,0,10,25,17,-28,6,6,20,41,14,-37,28,-14,-23,4,-27,-59,48,37,23,-18),
	(19,-62,-11,-3,-5,4,19,0,3,-27,-41,10,-60,-18,-38,39,59,-2,-26,-14,-9,-17,-53,8,-8,5,23,-27,-3,19,7,-4,31,-15,-4,37,10,10,7,11,-14,-26,20,0,32,-14,59,20,-3,41,9,21,3,-14,-14,-17,17,-14,19,14,-2,9,30,29,27,2,0,14,50,-28,20,-39,20,-4,0,33,17,2,-1,5,-7,17,3,25,-6,14,30,14,-16,25,-21,13,2,12,-20,-2,-12,-5,44,-1,17,21,6,1,-4,39,10,-17,27,6,-1,-49,20,8,23,5,-4,-37,41,3,-20,26,-22,-101,41,-4,14,14),
	(27,-23,-29,20,-19,30,4,-15,14,-36,10,-17,-21,20,-26,9,-6,24,-22,8,-13,-35,-67,12,12,29,7,10,27,-4,16,0,2,-25,-22,51,-16,23,25,-13,-39,0,18,2,14,-31,66,35,-16,37,-41,15,-30,-3,11,17,31,16,-6,-22,-8,20,-9,24,38,2,-1,23,33,-44,15,-5,0,3,4,11,12,11,-6,-9,11,-7,8,53,33,-7,16,-16,-11,14,-19,36,-8,0,8,41,-24,16,7,8,9,3,25,17,27,4,24,-17,11,2,15,-14,6,11,12,11,29,-18,46,-10,-29,11,0,-109,25,-27,15,-9),
	(32,-4,-24,3,-24,9,-9,23,34,-17,-12,-3,-1,21,-20,1,0,15,-2,-23,-18,-34,-64,29,0,25,24,20,33,-2,0,8,9,-11,36,46,-1,43,19,6,-10,45,20,7,20,1,58,9,0,-5,-21,21,-38,1,27,29,23,-6,-30,-22,-4,31,-23,18,50,-3,16,29,30,-44,29,30,-6,15,18,17,21,-1,9,10,-5,22,-11,38,21,-6,18,10,4,9,-19,0,-31,-25,0,7,0,23,-15,49,2,3,-5,40,33,-1,19,29,48,-41,-5,-24,23,20,10,32,8,8,25,21,2,-3,34,-48,12,-18,14,-5),
	(28,-18,0,7,10,28,25,15,11,-11,-8,-2,5,8,20,-34,-30,15,15,-30,4,-32,-27,32,-1,40,13,32,9,-2,5,22,-8,16,0,35,-15,14,18,25,-7,7,3,7,11,21,19,14,-9,24,5,0,-12,13,15,19,27,-7,-32,-22,11,7,-32,-6,35,-2,4,-9,24,-10,3,3,-10,14,22,-16,17,11,18,17,1,10,0,44,-3,19,-9,19,19,-9,26,21,-8,-40,-12,27,-26,43,-2,18,10,-14,-16,25,2,-13,18,16,18,-19,11,-38,31,14,-1,-10,17,-22,34,-10,1,10,39,4,22,0,-12,3),
	(29,-9,12,-7,18,10,-8,18,24,-15,-32,-26,7,25,29,-25,-7,-6,-3,-23,-10,-61,-23,21,-18,18,10,24,21,-41,-3,12,0,12,20,17,12,-7,30,14,-24,-16,14,18,7,29,-19,35,7,6,-9,-14,-17,-13,19,13,-2,-29,-38,15,0,5,-5,-7,46,-13,-8,-1,30,-13,24,-13,-18,21,9,-13,4,11,36,13,15,4,11,23,-22,38,13,21,17,-21,27,-27,-7,-41,3,9,-6,44,-31,17,28,-16,-18,-7,-15,-3,25,10,14,-7,16,-28,20,0,0,5,-16,-21,10,-19,4,7,25,-7,12,12,-9,29),
	(-4,1,1,3,0,26,0,2,30,-9,-37,-8,12,7,26,-47,17,-5,-4,-15,-11,-4,2,-17,-10,4,15,-15,5,-7,0,-8,10,18,-12,-20,-8,6,1,0,2,-39,-3,-11,19,3,-14,26,28,1,0,-16,-11,-14,12,48,-7,10,9,-14,0,17,-8,34,20,10,-6,-23,24,-20,9,1,-42,26,15,-10,17,11,12,11,19,12,8,45,-24,54,7,7,1,-30,22,-3,-16,-3,11,17,-3,21,-1,31,14,2,7,-23,-4,-13,42,5,21,29,18,-66,20,2,18,-1,-25,1,15,6,-13,-17,32,6,30,-11,-26,16),
	(0,0,11,1,-15,13,30,-29,-18,-2,-29,0,31,45,39,-26,-3,-16,-15,-20,3,16,-7,-6,-18,-26,0,6,-18,-24,-31,-14,34,21,-16,-45,-8,-32,-4,23,-7,-10,7,15,27,-6,12,11,13,0,24,-7,11,-1,-8,31,-16,12,28,3,-14,-5,-8,21,-35,26,-34,-8,-13,-22,0,-16,-33,15,-1,-8,9,10,3,14,-24,0,29,32,4,66,11,-1,26,6,-2,-26,-26,6,37,7,-16,17,26,-11,7,17,-15,-16,-20,11,20,22,0,48,25,-34,6,-16,-1,17,16,22,-22,14,-10,-17,1,-6,26,29,-23,7),
	(-29,3,16,-23,27,9,12,-28,-22,6,-21,-26,-13,3,32,-28,31,-31,1,0,-26,14,-30,10,-6,-27,-4,11,-4,-46,-20,2,22,17,-26,-40,9,-17,1,0,-11,17,18,-2,-7,3,33,-6,32,7,11,-8,6,0,-27,27,7,-8,20,-6,22,-12,-10,0,-89,23,-32,-17,10,-23,7,-6,-20,-3,-2,-2,-2,-14,13,-2,0,14,28,56,-18,47,19,-5,3,10,-28,-23,-17,-3,25,-19,-13,52,25,13,-9,17,-18,-44,-10,-24,-10,25,13,25,14,15,0,-14,-5,-1,14,-8,-23,20,4,-22,-26,-23,29,14,-8,6),
	(-19,19,-12,-8,3,2,29,-29,1,4,-17,-35,0,0,15,-27,10,-29,-21,-31,5,27,-20,8,10,-23,4,8,0,-53,-6,10,20,25,-22,-46,12,-14,-7,29,-14,6,-5,-9,9,20,2,1,24,11,11,-18,11,22,-27,12,-2,12,24,-7,18,2,-6,20,-94,14,-6,1,0,-23,-14,-37,-1,-7,-5,-24,16,7,24,-12,-9,30,21,20,-4,9,9,19,-14,29,9,10,-39,10,9,-17,-14,38,36,1,-1,-1,-1,-8,-35,-7,-6,12,-8,33,-10,56,-17,-11,8,5,-9,1,-2,20,0,0,-14,-43,-2,17,-28,2),
	(-63,3,1,-32,-17,8,28,-21,-11,15,-10,-12,-10,-36,30,-28,20,-38,-28,2,14,22,-12,26,17,6,0,-16,15,-49,-28,26,3,3,-8,-26,-20,-5,4,16,23,26,23,-26,-10,46,-15,11,-7,16,21,-3,0,28,0,-6,-36,23,20,-12,38,-4,7,5,-16,10,-38,12,23,0,2,-13,-8,-31,4,-13,-22,-5,26,15,13,-20,2,31,-13,11,13,21,7,36,15,17,-2,11,-12,-42,6,28,9,-7,-9,22,38,-39,-33,-10,-10,17,-4,-3,-28,33,12,-10,-18,9,8,9,-12,26,6,-15,9,-6,3,27,-11,7),
	(-58,26,7,-36,13,-2,30,-35,7,6,-3,-8,-39,-54,18,-5,21,-34,-22,3,9,-3,-8,0,7,-12,-12,-2,14,-40,-18,18,-30,8,-13,-29,-1,-9,-28,0,13,8,9,-14,-9,42,10,26,0,-4,19,-13,-2,10,-1,-3,-53,-9,22,-5,17,2,-29,-1,-32,-1,-28,-4,-5,-9,-20,-64,-42,-14,3,25,3,13,8,4,-6,3,15,12,-35,-3,29,13,-20,28,17,6,32,18,0,-21,17,29,-45,-21,27,30,5,-56,18,24,-23,-2,-32,24,-15,50,-17,-10,-13,29,9,6,-2,-10,-15,18,12,-12,37,-3,-10,-17),
	(-43,47,-4,-44,-10,-17,0,-21,-2,43,-18,19,-27,-26,16,11,22,-35,-11,10,24,25,0,3,39,3,6,-22,26,0,-15,20,-29,0,10,-28,-1,-7,-49,5,28,-26,43,0,-48,-10,40,3,19,-13,0,3,6,1,-18,-26,-36,10,-7,-20,11,-6,-37,-10,-7,24,-31,22,52,26,-25,-27,-44,22,-6,28,0,-48,-7,-1,-3,-30,5,-31,-27,2,17,23,-30,10,-17,-15,50,26,-11,-63,30,0,-72,-27,-7,23,2,-34,25,3,-42,24,-40,-11,-34,9,-9,-2,-9,5,14,2,-25,-5,-36,14,3,24,34,4,2,-21),
	(-36,22,10,-35,0,-5,-10,-19,-7,66,-19,70,-16,-41,-46,8,35,-34,4,-1,18,21,24,4,18,-7,-29,-35,15,23,3,-4,-39,9,-9,-16,26,9,-21,8,32,-14,37,15,-26,-7,15,-4,7,-36,28,23,-3,-7,-10,-7,-46,-7,-2,4,-31,-20,-29,-29,8,-16,-41,27,46,19,-11,0,-37,-8,-8,36,-12,-39,-36,34,-22,-49,16,0,11,-13,10,5,-16,-13,7,-9,34,16,-28,-37,39,-6,-23,-80,29,15,-51,-17,-9,19,-13,2,-42,-9,-54,12,-2,3,-9,20,17,-6,-15,2,-9,46,16,-50,28,-24,9,-7),
	(-18,5,0,10,-10,8,44,20,24,14,16,12,-46,-44,-29,44,21,4,-4,6,8,-20,15,-5,-39,3,-13,-14,-8,13,-18,-2,-14,-22,-26,15,-11,7,-23,-7,-11,-8,15,25,-7,-11,9,8,-43,-6,37,17,-10,-35,33,17,-12,-17,-23,-1,-31,8,17,7,-21,-43,-43,3,26,-38,26,-2,-59,25,18,20,5,-38,-18,57,-24,-11,56,-4,-34,-34,-11,0,-51,-5,-16,-13,-5,9,18,-20,57,-25,-39,-14,49,6,-47,-5,9,31,13,-12,3,-16,-20,-1,-6,2,-10,-12,-8,-24,-29,-17,-29,49,23,28,33,12,0,10),
	(37,-16,-32,16,-24,32,37,-17,20,-8,32,-55,14,-2,-9,15,12,12,-15,9,51,-1,26,-42,-31,60,-55,6,-15,-29,47,-27,29,-22,83,-16,27,30,-19,4,-8,-38,54,60,-34,-33,32,50,-52,-21,5,31,-48,46,26,47,-38,30,-58,13,-23,20,20,-10,-39,-31,-49,-7,44,-1,25,-12,-32,29,-18,45,65,10,-24,54,-31,27,55,-11,16,-28,11,9,-46,-24,-36,-27,-47,41,-22,-13,-18,26,-27,-27,50,-21,-18,27,-5,24,-25,-49,-60,-40,-2,13,-26,-30,18,62,8,26,-46,4,32,54,46,4,23,-17,44,-15),
	(22,-25,4,-1,-7,25,26,16,23,11,12,-27,7,0,-20,-9,3,28,-7,28,17,-19,0,-25,-30,21,-4,-1,-1,9,-2,-13,-5,-3,29,-1,-4,14,7,10,-24,-14,30,4,-32,9,2,-9,-27,-10,7,3,6,25,2,8,-22,-19,3,3,-14,16,-12,0,16,-30,14,-15,24,6,5,-4,-15,2,-11,-1,25,16,-28,31,5,7,18,-28,9,3,-10,11,-18,-11,1,8,7,35,19,-3,-13,18,-28,-16,3,-29,-2,9,-11,7,5,0,5,-21,-9,-7,-21,-11,7,26,-3,-3,1,-15,21,-5,1,-3,23,11,15,7),
	(7,-15,14,0,8,-18,-22,2,-9,-17,9,7,-5,15,-27,-10,13,12,-3,-5,4,-10,8,-1,0,-2,-19,3,-5,4,4,-8,-8,18,-14,13,-9,10,-18,22,10,-5,-7,-22,-19,-13,-3,-10,22,-21,-8,11,7,19,0,11,-1,-4,12,-3,4,-1,-13,-24,-25,17,9,0,-7,7,-16,-8,-14,9,-12,-18,5,-11,7,-7,16,0,12,-15,-6,8,0,18,-7,7,12,-21,-21,15,9,-10,3,-7,22,4,15,15,-24,9,-11,17,2,1,10,13,1,13,9,-4,1,-25,10,-13,-4,0,0,-4,15,10,-12,-6,-2,-17),
	(-11,-9,-5,7,5,2,-16,-6,13,6,5,0,6,-2,12,2,32,5,12,20,16,7,20,3,-14,-11,-3,-20,20,8,4,19,24,10,-1,24,-17,9,20,7,16,-28,-3,-3,15,3,-9,0,27,6,-16,12,-1,-5,0,4,17,24,-1,19,4,-22,9,-8,-16,-6,2,-5,6,-21,5,25,-16,19,-8,7,-14,3,-15,-7,20,2,-25,28,-6,2,-1,0,2,-1,-20,25,-6,10,-1,-8,-6,15,28,1,-15,0,20,-8,10,11,26,27,32,-11,-14,-11,-2,-1,24,5,8,-11,8,18,-27,-22,10,-11,0,-9,-13,16),
	(22,18,3,10,27,18,-57,27,-8,32,15,9,4,0,-18,-20,34,0,15,11,4,26,56,17,-23,-14,41,-51,20,24,-8,17,-25,-10,-8,34,-27,52,7,42,-6,4,5,32,5,8,-8,23,5,7,0,23,-3,-46,-2,-18,-1,10,-38,12,7,0,-41,26,25,-47,-25,22,-7,31,-9,23,-23,-24,29,-4,-22,-13,-6,-6,21,-14,30,13,26,2,25,53,15,-16,34,-5,-33,-2,-35,-3,-3,-36,-4,11,7,36,-23,12,-15,13,-33,-40,9,-12,-38,-48,51,24,5,-24,-31,15,-4,31,21,15,-9,55,4,-50,-10,1),
	(-23,-19,15,20,-2,42,10,-8,8,8,-20,-31,-7,-9,32,-4,41,1,27,4,-12,6,-21,-6,-41,17,11,13,2,-17,14,-6,-9,-45,23,-1,-1,-8,0,14,-34,13,44,-6,2,-2,-20,36,-21,-21,4,21,-14,-25,41,74,-29,-2,-9,-15,-33,42,26,4,-20,-5,-11,-42,-35,5,-12,-21,-11,18,0,-5,26,-11,36,20,-18,-16,46,-11,-5,-14,54,14,0,37,0,-32,7,-32,-4,-17,6,31,-29,4,19,-7,-44,-45,-6,-7,25,-30,-8,-17,-7,18,-10,12,60,-19,-13,-15,-19,3,-30,18,11,32,16,-55,-20,-18),
	(14,9,8,16,48,4,-33,21,-28,5,-59,7,-47,1,9,-28,9,2,-7,-12,-11,-27,8,-24,21,-10,-7,17,-2,-17,-7,-42,34,-47,-23,-63,-3,-7,-40,22,18,-14,-12,-27,14,-14,-40,19,-3,2,-28,33,-2,-34,-4,30,-14,1,0,-6,-4,61,15,-4,10,10,-4,-21,-33,-18,-29,-11,11,7,-36,-39,-1,9,-9,-27,-6,33,25,32,-6,-1,9,4,-18,22,5,12,1,8,16,-15,0,12,22,-4,21,-4,21,-40,-29,-9,-18,-51,0,3,-7,28,-16,-8,9,16,-20,16,-34,4,-24,8,14,-5,10,-43,-18,3),
	(38,42,23,15,14,21,-16,0,-50,14,-61,-15,-48,5,11,-21,18,-30,-42,-14,13,4,15,-25,12,-8,23,10,14,-31,-11,-25,-14,-13,-15,-55,-17,-26,-27,34,7,-14,-21,-50,15,-22,-20,11,-17,-4,33,35,2,-32,-40,12,-33,29,18,16,36,84,-6,-2,-15,12,9,-4,-17,10,1,-18,48,-5,-33,-14,7,-13,-23,16,-3,4,3,-25,-10,-21,0,-9,-16,5,-14,-11,16,21,-11,-7,-15,0,1,-7,20,4,0,-25,-26,35,-2,0,-40,-8,-37,20,13,-28,-20,48,10,-2,-25,-39,-42,-31,-8,-6,11,-3,-23,-7),
	(17,43,37,21,-12,16,16,-12,-43,47,-81,-9,-29,-6,13,19,47,9,-28,-23,14,0,-3,-34,-13,-5,4,-21,-10,-8,25,3,-25,-43,-26,-20,14,-5,-33,12,-29,6,-31,-54,31,7,-14,20,15,-34,10,34,-6,-19,-62,21,-41,0,17,3,-7,73,0,-10,-35,8,36,6,-42,1,23,-14,49,0,12,-12,-3,13,13,-4,-14,-1,12,-15,-6,-6,15,-10,-32,-2,3,-22,-14,-2,-8,-17,4,13,-35,-1,11,-14,1,-16,-32,14,-14,0,-45,10,-3,18,14,-11,-6,26,-4,-49,-48,-58,-55,-3,-19,-8,-6,-18,-35,-7),
	(38,58,31,0,15,17,2,15,-32,33,-72,13,-31,21,19,0,12,-1,-34,7,-21,31,29,-16,-2,-1,9,12,-7,-36,-18,-23,-30,-16,-30,-34,3,-23,-33,3,-10,-6,-9,-26,22,0,1,44,10,4,10,16,15,-43,-46,10,-54,5,6,7,-2,18,14,13,-89,11,29,-6,15,15,-18,-10,34,-22,-10,-22,-12,-19,26,32,26,-9,23,-16,-9,6,-4,-22,17,3,30,6,4,34,3,-20,-3,-11,-20,10,19,4,-1,-18,-5,8,32,-13,0,10,-11,-22,12,-7,10,13,6,-64,-36,-28,-28,-30,-16,5,20,-10,-7,-19),
	(35,43,38,13,10,21,22,12,-38,24,-96,12,-7,51,0,27,-1,3,-55,-10,-9,18,24,-19,0,8,-5,-8,14,-3,-10,0,-17,0,-4,-29,-20,-20,-12,-9,-52,8,-37,9,17,25,-46,55,-16,18,36,12,-22,-13,-54,34,-27,1,29,-4,-9,10,36,26,-43,7,-6,-12,45,14,0,-8,2,13,-2,-33,-2,0,17,27,9,-5,32,-14,5,22,-6,-12,5,31,4,1,15,38,-5,-1,-1,5,-22,9,32,9,-2,-8,-23,33,34,-24,10,18,17,-3,32,-11,21,-4,6,-61,1,-19,-24,2,-26,-5,3,10,-16,-15),
	(-8,-5,65,0,34,17,13,22,-12,-15,-106,27,-42,7,-2,0,18,2,-55,9,18,7,-7,-15,12,-11,-9,-11,11,-6,-16,-14,-32,-3,6,-25,-13,-28,7,-40,-28,-13,-13,-2,8,16,-55,29,9,2,58,1,25,-3,-34,0,2,-11,3,13,-25,13,31,1,-4,11,-28,5,30,29,13,5,-30,-13,-29,2,21,-12,5,-8,-1,-6,36,-4,-19,22,29,-6,31,10,41,-14,21,0,-6,-25,-30,-22,-16,-16,20,-7,4,-7,-21,9,33,-26,-5,1,-15,-18,3,-49,27,9,-13,-34,-12,1,-17,18,-20,-21,32,-1,10,-5),
	(10,-6,39,-23,-8,2,16,-11,-41,10,-68,22,-25,15,9,28,40,4,-50,11,0,-25,-24,2,27,8,15,-22,-18,33,-28,2,-3,-5,-15,-15,6,-51,53,-8,-37,-1,7,21,3,6,-21,27,10,2,49,-11,16,8,-35,11,2,-23,4,9,-23,20,32,15,22,31,1,6,70,9,-24,-24,-16,-20,-25,7,3,-30,28,0,0,13,-4,2,-24,18,30,0,30,10,16,-4,14,-2,-19,19,-63,5,-30,-35,37,26,-17,-13,-7,16,18,-6,15,38,-10,-35,-5,-4,30,2,5,-20,28,-14,-12,20,-27,-68,31,10,11,-16),
	(6,-52,35,-4,9,25,7,-25,11,-57,-10,48,-23,-5,7,20,30,9,-39,-1,-15,-26,-34,-32,10,11,-2,-7,-2,0,-9,5,7,-16,-18,-17,-4,-36,30,4,-9,-6,43,17,26,-15,52,-18,-4,-12,14,6,16,-19,-26,-6,6,-23,-13,-16,6,-2,6,29,12,10,-14,-2,53,-22,3,-25,-10,1,-15,28,25,0,-9,24,-7,0,9,24,-15,35,17,-15,0,16,24,5,19,33,-17,0,-65,32,-2,1,33,9,-18,0,0,29,27,2,29,33,-6,-22,25,-16,37,12,30,-13,29,-20,-28,41,-14,-121,40,3,34,-15),
	(0,-56,34,21,1,21,10,-37,-16,-30,28,31,-12,-17,-27,17,13,-4,-14,-11,10,-19,-23,-13,-12,-2,18,-20,6,26,-2,-22,-7,11,3,24,4,-2,32,-16,-25,14,20,13,20,-13,68,-17,9,9,-15,12,7,5,-12,-10,9,-22,-22,-12,-16,0,-19,36,51,2,15,40,43,-43,21,-7,26,-23,-38,24,-6,-23,-16,11,23,24,12,24,2,19,5,11,1,-3,-24,0,3,-13,-1,4,-45,-12,32,17,40,0,9,31,3,38,2,-4,13,-9,-10,-46,45,22,32,35,1,-4,47,-19,-23,11,-6,-153,42,-14,9,-10),
	(9,-25,-15,1,-2,25,-5,-16,33,-69,27,-6,2,14,-24,12,28,10,-4,2,-2,-17,-23,40,-25,28,7,18,13,-17,0,3,-16,0,19,11,-16,3,31,7,-32,15,26,25,29,-28,82,11,0,8,-51,-3,-28,10,-12,1,-12,-24,-7,7,-9,-14,-13,25,19,-36,-10,34,36,-31,44,21,-11,-15,13,-18,14,18,-15,7,-10,12,20,49,13,-39,12,-9,-11,26,-17,20,14,-4,-12,6,-40,10,16,9,51,22,3,24,39,10,16,18,24,-43,5,-2,34,-1,56,4,3,-14,22,-8,-15,7,27,-101,20,0,5,-7),
	(41,-7,-20,14,7,34,14,0,50,-10,37,21,-1,8,-39,12,-14,18,21,-17,3,-25,-35,35,-33,15,20,-4,21,-21,-11,25,19,-6,31,30,-16,43,-10,-14,-28,47,20,1,8,-17,51,32,-9,-7,-37,-1,-15,14,2,0,-21,-18,-24,-15,-32,-10,-35,-9,20,-17,28,-2,51,-22,50,42,-40,9,-2,-10,-4,4,1,26,-3,3,11,37,11,-32,-4,-13,-6,0,10,-9,10,3,-14,19,-26,7,-16,48,18,9,-1,33,33,3,0,15,22,-27,10,-12,9,29,34,3,14,-32,23,6,-32,3,-1,-25,10,-39,-14,-11),
	(11,-30,2,-5,-8,3,33,44,34,-19,-25,-15,12,18,2,-26,7,-4,13,-17,-29,-58,-18,18,-13,32,27,4,41,-25,-7,2,-12,-21,25,28,-4,4,-8,9,-5,-11,-12,-8,1,10,8,43,-9,-6,-18,-7,-28,3,44,18,2,9,-20,-2,-15,-1,5,2,9,-8,10,-8,23,-10,0,18,-31,22,-10,-12,-11,8,7,29,-1,11,14,24,2,9,6,5,29,14,14,-9,-4,-42,4,11,-25,31,-30,37,29,1,-17,-24,-3,-12,13,48,29,2,-12,-37,33,6,50,20,15,-20,9,-21,-18,-31,23,-8,26,-4,-12,3),
	(-1,-26,5,7,31,37,-1,49,14,-24,-43,-26,-4,-6,27,-12,-4,-16,-17,-3,-4,-50,-20,1,-13,-2,16,18,4,5,-8,18,-15,-9,11,-1,16,14,-6,-10,-18,-36,-2,23,8,31,-25,42,-18,-21,23,2,-19,-18,0,19,21,5,-33,16,-14,15,0,22,55,-1,1,5,12,-34,22,-24,-35,41,4,5,20,-2,10,7,-10,-10,37,19,-30,27,3,17,19,-12,26,-13,-18,-7,16,11,8,3,-3,-3,9,-16,-20,-3,-29,14,11,20,47,1,7,-57,4,16,0,19,11,0,9,-1,-31,-7,24,8,44,-20,-4,34),
	(4,-12,34,6,-3,14,24,18,-5,-30,-53,-8,1,20,43,-33,15,3,0,-1,-5,-2,-7,-9,3,-1,21,14,-14,-9,6,8,7,4,-5,-33,28,-17,6,-11,-38,-21,-4,-15,30,36,-17,14,18,-8,22,5,-2,0,18,21,30,4,36,-22,14,21,-7,-9,-9,39,-34,-27,-8,-7,-11,9,0,34,-4,-1,9,-18,20,-2,13,-5,30,14,-19,64,9,1,-9,2,23,-9,-29,10,44,-5,3,31,18,1,-7,18,-22,-38,-13,-9,18,-1,40,52,19,-35,13,-20,15,-14,-9,-7,-21,-2,-9,-22,22,16,20,0,1,25),
	(-4,-13,16,-21,-19,5,20,-6,-5,-23,-34,-12,1,16,17,-36,7,-24,-6,-18,18,7,-1,-7,17,-8,24,0,9,11,5,9,21,21,-30,-31,23,-24,24,17,-19,14,9,-23,-6,1,-5,-2,23,-6,22,10,-8,-5,3,11,34,14,26,-17,11,-11,-21,11,-41,21,-23,-4,12,6,-1,-10,6,5,21,8,-4,-2,10,27,-17,-4,26,30,-6,44,48,-25,0,2,5,7,-16,-16,37,3,-3,61,49,-27,-15,4,-17,-34,-16,-16,1,26,25,23,19,11,-21,8,-13,24,18,4,-9,-7,-4,1,-22,-22,16,2,-9,11),
	(-22,-14,-12,-29,5,-7,29,-25,0,-14,-60,-11,-23,-5,34,-50,13,-14,0,-12,1,19,-6,-25,-22,-16,12,-10,35,-40,-16,0,-4,24,-7,-17,-17,-4,-5,21,9,-12,-2,-28,26,-16,30,-19,-1,12,27,-4,-8,2,-39,41,3,23,3,7,3,7,1,6,-100,24,-22,-14,14,-35,12,-3,1,0,15,15,1,-18,42,31,-18,17,15,21,-29,40,12,22,0,-6,4,-10,-14,-10,0,-6,4,47,34,9,15,9,-17,-24,2,-3,-2,23,-20,12,-6,20,-11,8,-16,-11,-1,12,-34,-9,-13,-10,-9,-11,26,15,-16,11),
	(-34,7,0,-13,18,-33,39,25,-25,-11,-27,-15,-28,-11,47,-23,8,-11,-21,-36,5,41,13,-24,12,8,-32,-19,2,-24,-2,19,18,11,-21,-15,5,1,0,32,-1,-14,25,-27,8,6,-20,-11,30,24,10,3,17,0,-27,11,-11,19,11,-3,25,-5,-46,-4,-40,-4,-18,-14,19,-17,8,-18,29,-3,0,28,-16,-13,36,4,-23,2,15,20,-5,13,16,16,14,28,1,22,-22,28,-9,-6,0,31,26,11,3,-20,0,-25,-35,-19,-6,23,-8,9,-9,39,20,27,-8,19,0,-23,0,28,7,-2,-37,3,15,8,-15,-14),
	(-17,22,23,-23,-7,-6,32,-23,3,18,-32,4,-25,-6,17,9,16,-26,-15,12,4,9,0,-12,-8,-7,8,-18,23,-26,-34,15,-11,2,10,-19,-9,17,-2,33,21,0,12,-32,-26,16,-18,-12,2,-5,32,-1,15,21,-9,-14,-23,-9,-1,-19,6,-15,-4,0,9,-13,-39,-10,33,-12,-29,-21,-26,0,31,14,-11,23,13,-9,-4,-35,24,26,-26,-13,16,25,5,27,-17,-10,-2,7,1,-36,15,42,21,-12,3,4,-1,-51,0,7,-28,7,-35,19,-18,10,-9,24,-10,19,0,-13,-28,21,21,-1,-6,-52,13,24,-6,-24),
	(-54,29,15,-4,19,1,3,-19,19,2,-41,2,-50,-24,36,-18,-1,-24,-13,5,-10,9,0,-4,-24,2,-18,-21,12,-31,-21,17,9,-11,13,-13,-9,3,-40,32,13,18,1,-44,-17,47,23,7,14,7,26,-26,-6,8,6,13,-6,21,16,10,0,-17,-16,19,7,0,-52,18,47,9,-22,-44,-37,23,4,48,-26,-12,20,35,6,-39,20,-30,-32,8,30,32,-4,48,6,-1,20,4,-7,-23,18,25,-9,12,-5,-13,26,-32,-33,5,1,27,-49,4,-6,2,7,25,-20,11,18,2,-32,36,-22,-15,-27,-28,11,0,-17,-7),
	(-10,19,24,-51,6,-13,-3,-7,-5,6,-18,53,-43,-51,10,-9,18,-20,5,8,10,33,17,-25,15,-14,7,-2,10,-11,-15,-5,6,-23,13,-31,-2,-14,-51,20,43,-16,10,-15,-22,17,21,-11,23,-12,17,10,23,-7,22,-7,-35,3,0,18,17,-19,-2,-11,-9,13,-34,2,54,28,-18,-42,-31,12,4,31,-20,-26,-7,0,0,-52,-1,-50,2,6,43,28,0,16,17,-3,37,11,-12,-33,33,-12,-38,13,-15,6,0,-39,-7,24,-23,12,-28,-25,-27,-17,10,25,-18,14,17,-19,-25,21,-38,-8,-9,-47,43,23,18,14),
	(-6,19,-5,-12,0,-16,7,-1,-6,41,9,36,1,-35,-49,48,-6,-15,-16,25,48,-14,8,-17,6,-11,-23,-16,-12,22,9,-5,14,-22,-16,10,9,-8,-27,0,28,-4,37,1,0,-33,47,8,-19,-43,52,18,0,-32,5,-26,-28,19,-28,16,-2,0,-3,-18,-5,-5,-54,17,52,2,11,-22,-33,14,-6,37,-23,-28,-57,30,-14,-43,13,-25,8,-39,24,34,-53,-17,-4,-1,3,27,2,-5,48,11,-26,-30,14,-16,-19,-25,0,34,-17,-10,-38,-17,-31,-2,4,-13,3,1,3,36,-23,21,-18,14,-16,-37,23,-4,52,-27),
	(28,38,-9,-7,4,40,25,21,14,-12,-2,19,-24,-74,-10,30,-15,11,-40,-8,2,-24,12,6,-3,13,-47,-24,-13,-18,-3,10,16,-17,1,6,7,-11,-52,-23,-19,-19,57,45,4,-34,17,46,-35,-22,2,-7,-3,-54,11,0,0,-11,-18,9,-52,-2,-4,13,-11,-23,-15,45,-15,-30,17,-36,-65,13,3,12,39,-10,-22,20,-24,13,60,-50,-10,-41,-33,12,2,-74,-8,-21,13,25,-14,-3,49,8,-30,-5,67,-10,-41,-12,-21,38,-24,-10,-24,3,-30,-27,26,-13,-72,1,29,7,-40,-10,3,85,15,17,33,3,31,1),
	(-4,-23,-12,7,21,56,18,-5,23,-63,20,-25,16,0,-16,-4,18,-24,-51,46,4,-18,10,-40,-29,9,-34,0,17,1,36,-26,-1,-48,9,-10,0,43,-22,29,-26,-14,-9,-9,1,-9,-21,24,-25,-6,-2,29,-66,-2,43,46,-16,15,-35,15,-21,19,-2,7,-20,-50,-29,-40,20,-24,20,26,-34,21,-34,11,48,14,10,46,-15,24,71,4,18,-29,31,42,-33,-28,-28,-32,-29,-2,0,24,36,31,-34,28,39,-15,-23,2,-14,28,4,-39,2,-9,-10,30,-8,-8,10,-7,-42,21,-5,36,5,34,5,10,26,-45,-18,3),
	(43,-20,-33,14,-18,41,9,-3,-1,-29,10,-8,12,-20,-25,19,42,21,-13,38,39,-4,7,-3,-37,23,14,18,19,6,16,7,6,-34,15,-12,9,5,-13,-14,0,-20,44,41,-3,-33,-13,34,-20,-27,0,32,-40,27,8,35,-19,20,-49,17,-12,27,32,13,0,-28,-1,-19,14,-9,31,12,-6,24,0,25,10,16,-9,3,5,-4,37,-7,4,-35,-13,22,-3,-11,-10,-4,-15,26,-34,-22,23,36,-32,-11,15,-28,-21,12,-11,44,-31,0,10,-19,-10,34,8,-3,19,-4,-18,19,-5,-1,8,25,9,21,47,-11,30,-10),
	(7,15,1,6,-15,5,-15,-19,16,14,0,-14,12,-13,12,-5,5,-1,9,-14,-1,3,-13,-20,17,15,3,-16,20,11,-1,9,17,-12,-17,15,13,13,2,-7,0,-11,-15,-14,-3,-17,2,0,14,-7,-8,8,8,-19,9,12,-18,3,6,11,18,7,-2,-10,-13,-7,9,-6,0,11,9,0,13,11,-22,17,8,-11,-16,7,11,17,14,-13,17,-16,-12,-5,-1,-7,11,-15,-7,-20,4,16,-9,-6,17,-13,-18,-1,-12,-16,0,-11,-14,10,19,7,-9,-9,17,-15,-12,-18,2,14,8,-11,10,1,0,12,0,-11,1,13),
	(0,1,11,15,6,17,-15,-8,3,-9,4,-5,-12,-5,12,-31,4,-9,10,9,-24,-15,12,-35,-19,18,5,20,26,27,-35,4,19,-10,-30,6,-14,26,4,30,16,-30,21,18,15,27,-1,-24,15,9,25,-9,7,12,15,-4,-6,31,-16,14,-6,19,2,29,3,-39,-33,-12,-1,-6,10,30,-16,22,33,-10,0,31,-6,24,23,10,-20,31,22,-27,-28,31,11,13,7,-7,17,5,-3,21,7,6,19,1,-29,-11,6,-2,-3,6,22,19,0,-25,-6,-21,19,33,-1,21,27,-3,7,11,-1,-7,-21,-9,-17,-21,-5,35),
	(14,29,-21,-13,4,0,-33,45,25,-9,12,33,-9,4,-26,-17,31,-3,4,9,-21,-13,37,3,-14,-4,7,-11,33,19,9,11,17,15,-4,8,-31,34,22,0,32,-5,-1,11,26,-9,-5,-9,5,-9,15,28,-6,0,10,-29,0,0,-22,6,20,13,-2,21,33,-48,-18,7,-1,-8,26,23,-11,19,37,0,-9,-4,-29,25,17,-17,16,-9,18,11,-7,36,2,-9,-10,-5,-57,-14,-12,-12,-19,-22,-4,25,6,-10,10,24,14,1,12,-24,-13,-23,3,-12,17,17,26,9,21,5,27,29,-11,-18,-11,54,22,-22,2,0),
	(7,-2,-29,23,17,16,-25,-32,4,3,-55,-6,-21,0,-18,-5,51,26,33,15,-13,-5,-14,-12,-11,13,-5,0,22,15,52,-4,28,-10,24,-3,15,27,-26,1,-16,-13,24,0,19,-25,0,36,-17,-9,26,13,-16,-18,43,27,-40,-17,-59,-2,-26,50,17,4,-7,-35,-22,5,-24,-7,0,25,-28,4,-1,-5,-2,7,-21,28,-35,-9,7,-49,4,-23,31,18,-3,28,7,-7,-13,-6,0,-32,5,38,-11,-27,13,-18,-21,8,-17,-1,-40,-40,-26,-32,-5,-5,15,-10,27,-17,-10,26,-35,21,-19,-17,-2,22,27,-54,-26,-31),
	(-2,-4,-2,-3,11,4,-20,13,-29,2,-92,-47,-48,-29,26,-4,3,6,-16,36,13,2,6,-6,15,-2,-8,4,-1,21,-3,-4,61,-10,4,-64,1,-19,-38,16,3,-48,24,-27,0,-7,-6,4,-13,11,16,6,11,-11,7,18,-21,18,23,-3,15,52,-14,-14,4,7,43,-13,-36,8,6,2,45,0,-20,-71,-5,31,-5,-4,-10,17,19,15,6,-25,-12,9,-10,17,-26,-10,-18,6,23,9,10,5,52,9,-12,-34,27,-31,-18,20,-13,-20,-34,-21,-28,9,-5,23,13,4,22,-20,-8,4,-47,-23,28,-16,-10,-32,-9,13),
	(20,33,37,9,11,26,-11,-5,-24,29,-98,-29,-20,6,23,0,37,3,-28,-6,25,16,26,8,-2,17,-34,16,-2,-32,28,8,22,-39,-2,-46,-11,-14,-10,15,-14,-40,-5,-55,16,-30,-3,13,-1,-34,29,31,5,-54,-27,13,-30,23,-14,2,15,77,-6,-18,-21,7,23,-7,-32,-17,-14,0,60,-36,-14,-13,-7,4,3,11,-5,-10,3,-23,1,-22,-33,14,-23,-2,-6,7,3,32,-8,-19,0,13,24,7,29,-12,10,-27,-17,16,-33,-6,-30,18,-14,1,5,1,-23,18,5,-37,-15,-18,-35,-31,-16,-5,-14,-6,3,-38),
	(38,51,34,-8,-3,22,4,-30,-36,-11,-97,-18,21,10,40,8,2,1,-33,1,-12,37,2,10,15,1,-17,-25,-4,-44,4,-4,-10,-23,-34,-33,13,6,-24,0,-43,-16,-8,-58,-7,-28,7,28,-24,-3,1,35,10,-25,-29,19,-45,0,2,6,-9,47,26,-12,-33,13,36,-1,23,-2,-9,-8,19,0,-17,-58,34,-17,22,24,-20,-16,40,-21,-16,-11,-40,-12,-20,0,11,-15,-8,4,5,-47,-38,12,-18,10,6,5,-15,8,-2,21,-1,22,-42,8,11,-16,21,-15,11,15,13,-48,-43,-45,-12,-25,-22,8,23,-3,-12,-5),
	(18,56,11,-11,27,24,22,-3,-17,33,-108,-7,-7,0,14,-4,34,0,-69,23,8,53,27,8,-5,7,-19,-3,8,-33,8,-11,-8,-12,-26,-14,5,-19,-29,0,-21,-28,-14,-48,-6,11,-16,22,-18,11,15,5,28,-42,-68,2,-23,12,24,-5,-7,19,21,32,-56,16,0,0,49,13,-5,-7,32,29,-2,-32,8,-15,33,47,12,-18,39,0,-33,-3,-40,-2,-2,-16,27,-9,-22,5,-13,-25,-22,-9,-29,-22,26,-18,-7,-20,-6,26,-10,2,-29,34,0,-28,4,-25,7,-7,-10,-61,-42,-43,-13,-31,-27,-10,33,-20,-6,-1),
	(16,40,49,-5,-1,39,29,-9,-5,-7,-115,15,-31,72,10,16,15,-7,-54,1,16,28,5,25,10,-15,0,-37,38,6,11,-12,-25,0,-41,-48,1,-16,-10,-29,-33,2,-23,11,0,21,-32,56,14,12,51,4,0,-28,-46,34,-20,-24,35,-6,9,3,19,12,-42,42,0,-27,70,21,10,-21,2,-9,-28,-72,27,-12,17,30,29,-30,9,-3,-17,22,-38,-18,27,23,12,-20,5,19,-27,-6,-19,-4,-39,0,5,-9,7,-31,-24,1,12,-23,-33,22,11,0,2,-31,-10,23,9,-49,-44,-58,4,-13,-19,-64,22,-23,0,-15),
	(20,24,46,3,24,2,29,13,-1,13,-60,0,-28,39,-17,26,16,-10,-33,4,-12,-12,7,-12,1,3,-31,-3,23,-5,0,3,-16,-40,-29,-29,3,-26,10,-16,-47,-3,-15,3,20,10,-6,22,-21,1,41,12,31,-39,-68,-1,-42,-5,7,-3,-21,-7,15,22,-50,15,-18,9,72,-12,21,-21,-12,-16,-10,-51,26,8,23,12,2,-6,24,15,3,11,-14,-10,34,32,22,-9,4,17,-27,-25,-16,6,-61,-14,38,0,13,-1,11,39,21,-45,-6,14,21,-15,29,-13,18,21,3,-45,-42,-22,11,15,-47,-70,25,-16,23,-10),
	(22,-3,43,0,-20,6,15,-11,0,2,-22,49,-31,23,18,22,29,5,-11,7,27,-26,-13,10,5,35,-28,9,-11,17,12,-15,-28,6,-8,-41,13,-15,30,-37,-10,-3,37,13,24,-5,26,-7,-17,-12,38,14,6,-1,-45,-3,-12,-18,5,1,-25,13,21,31,6,29,-12,0,76,5,26,-6,-31,9,-53,-34,34,15,-7,6,14,-14,-3,22,-9,14,-34,-29,29,24,-4,-5,2,27,-9,30,-31,28,-41,-32,11,-23,27,15,-7,47,8,-13,24,2,-5,-25,33,-21,31,32,2,-32,0,-29,11,17,-25,-105,41,-11,24,-34),
	(33,-30,42,6,8,23,5,12,-9,-32,6,31,-40,25,-15,17,19,3,7,-18,24,-63,-25,-8,-15,15,10,4,10,8,18,-8,-5,21,17,-11,-16,-26,44,-38,-27,5,50,23,0,20,71,-32,1,-21,25,18,-19,-10,-39,14,-30,-5,6,-2,-7,0,11,30,23,-6,-10,35,55,-35,29,-13,-40,1,-29,-11,25,-24,-10,25,34,33,5,43,-10,12,-12,-8,44,15,3,16,11,5,-3,40,-36,13,8,-25,39,4,-9,9,27,12,-17,3,36,18,13,-6,41,-16,7,3,16,-41,0,-22,-17,46,10,-185,46,21,40,-11),
	(9,-41,29,-5,1,10,10,-20,-9,-46,47,25,12,7,-23,4,18,24,20,-13,-3,-25,-33,0,-8,34,28,9,21,7,-7,-5,18,-25,7,-9,-5,-14,43,15,-31,37,10,32,19,-21,79,-27,-24,0,-45,17,0,14,-45,9,15,-4,-14,1,-28,-20,-7,26,0,-23,-8,28,60,-30,23,0,-9,-7,-45,-10,8,8,-16,-6,1,30,19,23,-3,22,17,-32,0,17,-24,0,22,1,6,8,-72,19,1,-31,40,13,-11,0,23,8,9,9,9,-9,24,2,31,-16,25,-1,24,-17,42,-14,13,39,-10,-133,0,14,12,-18),
	(12,-37,-1,18,6,31,-15,-12,3,-49,59,13,0,13,-50,0,15,13,27,16,-16,-18,-8,9,-3,43,26,17,31,-2,18,-22,4,-5,28,4,-3,26,31,-17,-28,42,6,11,12,0,38,21,14,17,-78,-6,-8,3,-18,32,9,10,-38,-7,-34,5,-27,9,-6,-8,16,21,65,-16,24,33,9,5,-7,-22,9,16,-10,22,14,-12,30,33,15,-15,-30,-19,18,17,-22,-26,0,0,-16,17,-41,23,12,24,34,11,-11,-1,14,1,-2,17,33,-38,12,-9,39,-2,39,7,17,-24,44,10,-9,21,19,-45,16,-20,-6,7),
	(18,-20,12,-3,-8,24,30,1,22,-18,38,14,31,-8,-8,11,14,2,7,-15,-36,-5,-43,11,-18,30,-4,-23,50,4,-2,18,-6,10,22,-5,10,27,11,-5,-30,34,18,24,13,10,53,48,-14,-17,-24,0,-20,9,16,27,4,-28,-4,-11,-37,2,-29,13,3,-20,22,-17,12,-13,34,10,-14,-14,3,-9,-1,2,7,18,3,-13,19,25,15,-12,-2,6,17,12,6,-29,-20,-5,8,-16,-49,-11,-22,46,24,10,6,2,16,26,-5,25,43,-26,-5,-1,11,20,40,0,4,-2,21,-2,-14,2,41,28,25,5,-19,0),
	(26,-9,19,16,25,8,4,-1,5,-19,-30,2,3,8,24,-12,0,-11,-14,-18,-21,-43,-4,-1,7,20,20,-18,23,-11,0,1,-11,-21,8,-13,6,22,-1,9,-18,11,7,-14,15,12,18,54,22,19,-3,13,-31,1,13,4,3,-12,-22,-21,-25,4,5,-23,7,18,19,-11,21,-6,-15,10,0,-6,-17,-29,26,14,20,3,12,-23,57,18,-12,29,-13,-20,-12,3,40,-39,-4,-18,6,-9,-17,4,-26,-12,17,25,0,-19,-38,17,24,45,28,30,4,-40,16,20,58,-18,0,-3,13,-7,-17,3,31,62,29,-15,-12,-15),
	(-7,-69,11,-10,26,39,2,-4,0,-35,-8,-3,-3,3,18,-3,11,8,-4,11,-6,-28,-17,-12,-11,17,-22,-10,-1,0,-1,-16,0,-7,18,-21,6,-9,21,-24,-24,-6,-13,22,26,0,20,26,19,-14,-5,1,-29,-20,24,32,0,-19,-17,-5,-15,-2,-4,-9,3,25,20,-7,-10,-18,0,-13,-2,4,8,17,34,7,10,0,18,-14,69,-14,0,54,1,-14,14,15,20,-18,4,6,24,29,32,-16,5,-27,37,13,-9,0,-25,-9,38,8,36,50,31,-40,20,-14,39,15,-12,-23,20,-12,-15,-19,5,20,48,-11,11,4),
	(-11,-39,3,6,-11,-6,29,9,0,-1,-29,-46,-5,-10,47,0,25,-33,6,16,-21,14,-1,-22,-18,12,-17,-14,-25,-4,3,-27,13,-18,-25,-32,18,-7,31,25,-5,-38,18,-6,9,-1,-16,20,31,17,3,11,-11,-2,6,21,36,-6,29,16,9,16,17,0,-36,39,15,0,-14,-12,-11,-11,9,17,-6,4,17,-11,32,23,18,1,41,2,-34,39,27,-22,16,-17,21,-25,11,-12,50,6,7,45,8,-9,37,-6,7,-9,-17,16,26,18,6,46,22,-37,0,21,-3,2,1,-8,12,-16,-21,1,-15,2,53,5,-9,20),
	(-28,-2,3,-21,11,6,6,24,-23,7,-26,-33,0,-15,42,-31,33,-41,0,11,4,0,6,-22,-17,-12,-15,-20,25,12,-14,14,-1,18,-23,-22,-11,5,10,37,-11,-2,-14,2,26,11,11,-10,20,1,8,-1,-27,22,-11,22,11,11,-3,-13,18,9,-17,14,-60,30,-19,-3,22,-23,-7,8,11,18,28,0,17,5,32,28,0,3,49,17,-14,56,12,-1,-8,16,14,1,-17,15,11,-5,24,38,24,-7,-14,-12,-12,-32,2,-20,-11,9,9,26,-1,-3,21,11,-6,-12,-4,-2,8,-11,-3,-13,-39,-28,14,-17,-29,11),
	(-23,-22,3,-22,29,-22,21,-10,-19,-1,-24,-23,-1,-11,30,-14,24,-13,22,1,-18,19,-4,-31,8,-5,9,-37,14,-8,-17,3,13,-2,-36,-28,22,10,-2,38,-10,-1,20,-8,14,-13,22,-5,36,-13,20,-18,-15,9,-4,-10,5,7,7,18,-7,-8,-12,0,-85,-6,-46,13,21,-14,-9,19,-2,14,26,35,-7,-29,40,1,-30,-6,21,48,-3,50,20,0,4,12,7,-1,3,19,-11,-5,15,47,31,-5,1,-8,-11,-14,-9,-19,-32,-10,-24,11,-15,32,6,30,-13,0,25,15,-22,1,14,6,-50,-13,18,-3,-40,-14),
	(-27,11,18,-54,13,1,14,20,-9,5,-48,9,-2,-20,23,-1,3,-20,-3,-15,-21,20,-1,-10,-8,-17,-31,0,26,-26,13,-3,14,12,-15,-10,23,11,-23,40,4,2,13,-43,21,7,-1,-15,35,-15,11,-5,-12,16,12,-10,-20,14,15,-13,25,0,-3,-14,-12,-3,-29,0,-1,-38,-7,5,5,13,-1,21,0,-14,23,21,-26,19,47,-4,-18,-3,5,26,-17,14,5,-10,-24,4,-3,-35,19,25,28,-6,-21,-25,-24,-11,-33,-27,-23,6,-41,35,-17,12,-13,7,-23,-6,-9,-6,-28,20,11,-16,-18,-13,-1,19,-24,7),
	(-8,-5,-3,-26,8,13,2,3,-20,-10,-6,0,7,-24,0,25,20,-11,-7,26,6,38,5,-7,10,-4,-26,-16,20,-62,-13,-14,7,-6,-5,-8,13,4,-26,8,17,23,-3,-18,10,26,19,13,2,-20,30,0,12,3,11,1,-50,-16,7,-11,-12,2,18,-5,17,9,-59,-14,28,-9,-5,-28,-56,19,17,61,23,3,5,22,-10,-32,68,-35,-21,-7,-7,54,-11,17,1,-39,-8,19,-11,-63,4,17,8,-28,33,-42,-35,-29,-6,-6,-6,-18,-15,-3,-1,-7,-13,-5,-2,-23,-6,22,-56,5,20,6,-7,22,32,14,-14,-40),
	(3,41,-2,-35,-21,-11,-12,-17,18,7,-9,28,-23,-15,-5,24,-14,-10,-19,0,-6,8,-14,-25,-19,-1,6,9,10,-35,-29,6,-4,-24,-23,-12,31,11,-47,20,2,20,0,-20,1,18,15,-17,-3,-2,-1,-7,-3,13,14,7,-33,10,-22,13,1,-11,-18,-13,14,-3,-69,-1,40,4,14,-5,-41,32,-8,64,11,8,3,26,-23,0,18,-61,10,-15,14,33,7,21,-21,21,9,10,-21,-3,27,32,-15,12,0,-3,16,-34,-15,5,-9,17,-23,10,-1,-23,-1,29,-2,8,7,3,-38,23,-1,3,1,0,36,-7,13,-18),
	(-20,32,5,-6,2,9,-17,-5,-2,-5,-1,27,-4,-46,-25,22,-8,-18,-31,1,4,4,-4,-17,-6,-9,-4,14,16,-10,-14,-25,4,-44,-13,-3,-18,18,-73,-3,-8,-1,8,-26,13,-13,23,14,5,-17,22,-12,22,-26,14,-19,-39,-19,-19,-14,-20,-54,20,-30,11,-1,-83,17,45,4,-6,-19,-66,19,7,46,14,-10,-28,20,-21,-37,15,-67,14,-16,6,19,-19,17,1,16,9,6,10,-23,54,27,-70,-26,5,-9,-26,-7,-3,29,-12,-21,-40,-26,17,-62,11,37,3,-7,16,-13,-55,-4,-23,12,-3,7,19,6,12,5),
	(-19,28,0,-26,2,-2,-29,5,3,22,40,46,2,-50,-39,53,7,-3,-40,30,18,23,-3,4,-10,24,-26,0,29,-15,0,-1,-4,-39,-29,0,14,23,-71,32,28,-17,23,-12,0,-38,29,-9,3,-4,32,-3,-12,1,25,-24,-53,0,-5,5,-28,-4,0,-28,13,-40,-24,15,31,2,10,-7,-73,9,13,41,-13,-7,-45,3,-17,-33,30,-57,0,-56,12,28,0,30,-9,-4,7,-2,4,-14,9,-19,-22,-17,-24,-4,-28,7,21,45,-17,4,-37,-12,-40,-17,18,15,-12,6,1,19,-24,4,-16,-8,9,-11,24,-21,10,0),
	(43,25,-20,8,20,88,48,-1,-17,-21,47,5,-9,-62,-17,36,2,-9,-24,32,4,-30,-8,-40,-46,60,-9,10,-13,-7,30,-5,2,-22,34,-15,-6,20,-50,-28,-38,-8,56,42,0,-48,38,77,-54,-17,-11,-4,-42,-36,0,0,-31,-22,-71,0,-42,-43,15,-8,-35,-47,10,33,5,-25,59,-20,-22,-26,-1,57,67,0,-30,30,-29,18,50,-40,-32,-26,9,19,-20,-70,0,-32,21,46,-19,-9,12,21,-44,-27,70,2,-50,-15,0,36,-45,13,-56,-9,-59,-17,42,-63,-54,5,3,-5,-51,-40,50,93,13,-11,36,3,26,-28),
	(40,-26,2,7,6,68,43,-3,11,-57,33,-56,10,-13,-44,17,12,18,-36,35,12,2,4,-32,-65,35,-10,26,20,-25,24,-16,1,-46,63,9,53,52,-43,-38,-39,-30,8,28,0,-64,-4,52,-34,-25,-17,57,-43,-7,54,29,-28,0,-59,0,-49,18,33,-19,6,-56,-10,-18,42,-27,4,20,-10,15,-29,21,35,0,-12,51,-24,-2,73,9,-2,-35,15,3,-66,-44,-75,-41,-42,32,-7,-34,-29,10,-38,21,46,-42,-23,-8,12,29,4,-47,-26,-35,-3,20,-20,-38,1,40,-41,17,-48,-5,6,95,6,12,51,-41,15,15),
	(13,-40,-25,5,-24,6,22,30,25,-17,19,-43,34,-9,-35,35,15,0,-28,5,7,23,-6,-13,-12,32,-12,9,-13,-24,21,-10,37,-10,13,-23,25,19,-29,-38,-5,-17,25,39,7,-31,-19,-9,-37,-41,10,19,-27,6,35,-9,-12,38,-6,-1,-10,14,24,-22,-29,-16,18,-16,13,-27,45,24,0,39,-33,13,25,15,-61,0,-20,7,24,-48,0,-30,15,-17,-17,-31,-44,-29,-38,46,-2,6,40,2,-36,-2,22,-31,-10,-4,7,32,-20,-2,-30,-1,-14,22,-41,2,-22,25,-5,38,-5,32,39,21,45,18,21,-15,36,-42),
	(-7,-12,7,5,2,7,2,7,-17,14,10,-10,18,-5,3,4,11,7,-10,13,17,10,-18,8,19,15,0,17,15,-9,-11,-14,-17,-17,-12,17,-2,13,7,-6,-18,-7,18,-10,12,0,19,6,-10,-18,-16,11,-3,-8,18,-1,6,-8,-11,-2,-8,1,14,8,15,-7,-14,2,15,-5,18,10,8,7,-15,-11,-20,-15,-19,19,-2,10,-13,-2,8,3,3,14,7,-2,-19,15,-3,6,15,-9,-12,13,8,-10,-6,-16,6,18,-14,-8,0,14,-5,-12,-13,-8,19,-16,-13,4,12,8,5,-16,17,7,9,-11,14,-16,17,-7),
	(-28,-9,-1,-14,21,4,-21,6,13,-11,8,7,10,-2,-24,1,7,0,23,7,-10,-16,0,-28,-31,1,-18,6,5,31,-4,32,-5,-16,5,15,-33,33,26,25,2,-9,18,-11,-14,-13,-9,-34,-6,16,-4,4,-24,13,19,-12,10,9,7,-6,20,13,3,12,28,-6,-19,15,9,-19,14,8,22,19,11,-8,-30,-2,-2,-19,-19,-3,9,16,-2,-20,-21,25,-8,21,-25,-10,18,-16,-36,29,-5,-8,5,32,-17,2,16,3,-13,-29,23,7,13,-15,-23,-13,4,8,30,26,6,32,22,32,-15,6,5,-7,10,-17,-30,8),
	(1,14,15,8,16,22,-5,17,14,8,-37,29,-5,-26,4,-9,43,8,12,24,-49,-6,8,-3,-41,7,4,-10,38,2,-19,-2,9,-47,2,15,-9,28,-23,24,-22,-41,-8,-12,11,-18,28,25,-17,28,-8,28,-39,-6,0,37,0,14,-19,-11,1,25,28,8,15,-40,-36,-13,-17,1,8,13,-20,-15,4,27,-8,-21,-1,60,-16,-2,17,7,1,12,29,1,23,9,19,-14,-15,11,-25,-29,-15,-4,8,-13,-5,-15,-2,3,-18,16,-11,-27,-1,-6,-6,0,32,17,41,-9,3,12,-3,9,-28,-15,-6,31,45,-32,-12,9),
	(27,7,-24,7,0,11,-10,2,20,-17,-53,-2,7,-53,-37,-25,35,2,29,42,-25,-22,-45,-22,-21,34,-15,10,1,25,49,22,37,22,14,-39,-15,63,-44,26,4,0,-9,-10,37,-20,4,11,-3,-8,18,59,-28,-13,20,14,-35,9,-39,8,8,46,23,-21,-3,-26,3,13,-34,-7,23,43,-13,-18,38,-22,2,12,-26,0,-18,46,5,-12,29,-33,6,19,-22,3,-3,3,-5,-11,-44,-1,8,45,18,-12,10,-10,3,32,-20,7,-17,-31,-3,-38,-37,-6,37,6,59,-3,22,34,2,24,6,-6,3,-7,19,-18,-8,12),
	(15,-4,-42,0,25,8,-4,9,-16,6,-73,-45,-1,-32,20,12,34,7,-14,31,-10,29,15,-22,-17,17,0,10,9,19,3,-21,29,-5,-11,-29,10,23,-31,9,-16,-8,0,-13,-7,-9,39,18,-4,-2,46,40,10,-24,-13,-4,5,0,20,-14,0,44,3,-27,9,-31,-2,-5,-52,-12,3,13,20,-16,1,-35,20,-4,-22,24,-17,12,21,-10,30,-27,-43,19,-8,-4,-8,-3,6,13,-38,-17,-8,20,51,18,-11,-43,-19,-7,-26,-2,-46,-25,-21,3,-34,4,-4,5,20,-21,-22,-15,-18,-4,-24,-37,-3,-2,21,-13,-10,-18),
	(9,19,-11,4,-2,-7,-18,-14,-24,-15,-82,-10,-35,18,3,18,17,-7,-34,15,21,27,19,-35,28,-10,-15,-10,-12,-34,37,8,0,0,-9,-41,0,12,-38,-2,-31,-37,10,-64,-8,-14,4,-4,-12,-4,20,18,4,-46,-15,6,-19,12,-6,-21,2,23,-13,-35,18,-13,48,-19,11,22,-5,0,44,-36,5,-57,30,-7,2,13,-15,26,26,-7,-16,-13,-50,21,-29,-20,-9,-22,14,8,-40,-13,-31,10,21,16,-15,-32,-9,-6,16,15,-56,-13,-41,8,-28,0,-4,17,25,-6,-16,-36,-43,-33,-19,-13,-22,-27,14,-11,12,-20),
	(32,44,13,10,-2,28,8,-16,0,2,-96,-17,-2,-19,14,14,1,18,-34,9,22,33,15,-17,15,28,-26,-4,17,-60,26,-15,24,-9,-35,-30,5,28,-33,-2,-42,12,-4,-76,-3,-10,-22,21,-15,-38,5,8,17,-29,-28,35,-23,-5,-3,-16,4,23,14,-24,-62,4,30,-32,0,13,-4,-28,33,-20,12,-23,33,-15,7,-3,-18,11,31,-32,-8,-28,-93,-22,-10,-40,-9,8,9,10,-16,-33,-25,20,23,-20,30,-4,-21,-1,10,27,-42,-34,-71,-11,-20,-1,-6,5,-12,7,-33,-54,-38,-53,-8,0,-34,-54,-12,-25,-8,-4),
	(5,48,18,-16,-2,-3,31,-32,6,-3,-48,-50,-12,9,17,-14,5,-6,-45,-3,9,37,18,13,-22,21,-34,7,35,-24,8,-29,-14,-21,-50,5,6,-9,-47,-19,-53,-42,-53,-76,-4,19,1,41,-1,-11,29,6,-8,-24,-42,26,-25,16,-2,-18,23,13,9,7,-61,21,2,6,22,-18,-20,-46,14,21,4,-39,2,-24,6,38,12,4,33,15,-21,-13,-93,-23,-13,-15,11,-18,-28,10,-12,-47,-25,33,10,15,8,-34,-8,-17,-8,-3,9,-28,-74,-5,-13,-11,26,-1,-7,-1,3,-57,-33,-47,-15,-18,-36,-29,-15,2,-2,-27),
	(36,60,22,25,7,2,49,-27,5,13,-48,-12,0,20,20,12,34,-4,-34,13,15,18,8,-2,-15,15,-47,-1,-4,-27,14,-29,-32,0,-31,-21,10,-10,-35,-9,-72,-18,-35,-24,3,-9,-2,19,-16,22,37,-4,19,-15,-46,30,-15,-7,2,12,-25,-9,23,29,-26,-6,-1,14,58,-14,2,-12,-9,-13,0,-42,7,-1,11,25,3,10,24,0,-10,19,-76,-32,13,-8,15,6,-6,19,-6,-43,-23,22,-14,-13,42,-33,-11,11,-4,29,-3,-27,-49,16,11,-25,22,-4,-11,-1,26,-64,-49,-65,20,2,-51,-74,5,-29,25,-19),
	(32,38,24,0,-3,16,14,-31,14,-27,1,6,-15,59,-34,0,20,-9,-26,-24,-8,-17,16,11,-7,-1,-16,-2,-18,-11,-10,-24,-41,-42,10,-33,5,-2,-31,-21,-69,8,-27,29,23,0,-8,-12,-24,-12,68,17,12,-43,-34,-11,-26,-8,24,12,-16,13,23,21,-26,13,4,13,58,-18,1,-12,-26,-19,-26,-61,31,-20,34,26,-8,8,29,-1,-28,13,-89,-15,31,-11,22,-18,-11,8,-21,-37,-9,8,-25,-5,19,-17,-23,-12,36,44,-3,-29,-40,20,15,-15,5,-29,8,4,-15,-28,-22,-70,-1,30,-19,-100,29,-5,30,-19),
	(16,35,19,14,-9,12,28,7,12,-7,9,0,-6,36,-23,28,16,11,2,-20,16,-1,23,8,-5,16,-9,2,-44,-1,22,-19,-28,-21,8,-48,-12,-21,0,-40,-35,-1,22,23,-3,22,38,-43,-22,-13,35,-3,15,-28,-60,-8,-13,-13,-4,11,-2,9,12,21,-14,19,-1,9,28,-30,25,-22,-16,5,-42,-75,5,-3,-26,19,23,-20,23,20,-25,20,-49,-17,13,-11,5,0,-11,31,-13,-9,-29,15,-30,-15,23,2,6,-15,34,35,-6,-37,-28,15,0,-18,16,-43,-2,27,2,-52,-19,-45,3,60,11,-159,13,-1,27,-19),
	(37,7,27,6,-19,20,12,-19,20,-24,35,10,4,29,-29,0,23,-6,26,1,1,-19,13,30,-19,18,3,17,4,3,22,15,-7,9,26,-36,3,0,-2,-20,-27,-7,41,0,35,-4,76,-46,-13,-12,3,23,-7,-20,-55,10,-28,-17,-24,0,-25,0,13,24,-7,4,-26,6,30,-20,-8,-15,10,-23,-66,-63,33,-7,-15,6,18,0,-1,30,-4,-5,-66,-20,33,-16,-26,4,2,1,3,7,-58,-4,8,-31,32,-3,6,-15,28,23,6,31,-35,-4,15,-1,32,-35,36,20,1,-27,-16,-50,-11,55,11,-157,11,23,24,-33),
	(5,8,11,0,-6,20,-4,-27,12,-29,66,33,11,47,-76,-5,-2,8,25,-15,-2,-29,-4,18,-4,33,10,-3,-3,-38,-11,-3,14,-14,15,-33,-22,5,9,-30,-61,38,63,30,9,-2,44,-39,6,-17,-39,4,-29,-23,-24,26,5,-5,-21,-3,-23,-4,-7,15,-1,-11,-34,7,66,-10,20,9,-4,9,-64,-69,11,-18,-17,34,0,9,25,29,-12,-20,-81,-29,31,-13,-34,8,-12,-3,15,-4,-59,-1,-20,-12,38,21,-3,5,35,39,6,38,1,-17,6,0,0,-6,38,-16,-4,-23,-10,-16,7,31,12,-88,21,-7,26,-25),
	(-6,-29,-10,30,-26,23,-5,-29,24,-37,61,19,16,55,-44,-10,2,8,28,-10,-11,-28,0,11,-11,36,-6,11,14,-12,7,7,14,-3,38,-18,-8,33,17,-13,-85,34,40,-11,2,8,51,18,6,17,-63,6,-20,-1,-9,12,-16,-25,0,-12,-29,6,-19,4,30,-22,-5,-22,46,-2,15,5,3,-1,1,-45,17,-7,15,17,-15,8,31,42,10,-26,-90,-34,22,30,-17,-33,20,9,-5,10,-38,8,17,23,10,54,-19,10,11,17,-1,28,14,-18,0,-32,4,-7,45,-19,0,-25,34,-24,-2,-12,45,-3,34,0,-22,-15),
	(20,-23,10,12,-7,13,13,-38,22,-18,27,16,35,7,27,-5,-8,-19,34,-20,-15,-19,-13,21,-7,32,-6,-24,17,1,20,14,-32,-12,6,-13,0,8,9,2,-43,10,-10,25,2,50,14,46,3,10,-49,11,-1,3,-12,27,-1,-10,3,-16,-31,-20,-2,-16,12,-8,24,-1,11,-12,-9,23,3,9,-15,-39,5,4,34,12,10,-35,42,10,-23,12,-63,-8,19,7,55,-24,-16,0,-6,-22,-68,-23,13,9,-12,19,-11,-15,-7,14,1,25,0,8,10,-24,-11,-7,12,4,10,-17,0,-28,-29,-18,14,30,25,-14,-11,-13),
	(20,-36,35,-7,-4,9,-3,-30,-8,-23,-4,-15,-19,17,41,-27,4,8,13,4,6,-33,-10,-6,-14,14,-17,-9,2,3,10,-12,-15,0,16,-18,19,6,4,-6,-2,16,9,-2,-12,28,2,26,1,8,-17,6,-18,-8,27,31,12,-12,14,-21,-2,0,-4,-5,-17,14,42,-1,21,-17,-2,-14,18,10,-16,-16,15,14,-5,8,27,-10,39,7,-19,56,-12,-22,-9,2,61,-30,-12,-9,-8,36,-15,-11,-24,-10,37,31,3,-14,-17,16,14,41,23,46,10,-58,-13,-15,11,-15,-33,-24,27,-1,-20,-9,28,42,43,-20,-13,-9),
	(-33,-57,27,13,31,0,28,14,-8,-34,2,-42,-10,-10,59,0,13,11,15,-3,-27,-21,3,-30,2,5,0,15,-18,16,-23,13,4,5,8,-6,27,-12,8,5,-15,-38,6,5,17,14,30,31,-3,24,-24,17,-8,-12,16,13,38,0,26,-1,-11,-13,-21,6,-19,11,20,-1,15,18,-12,-8,9,0,-6,0,19,-4,15,2,-7,-19,72,5,-17,40,20,-6,-4,19,33,-21,15,-5,30,27,25,-16,8,-53,4,19,-3,-17,-22,13,-6,39,4,40,-3,-42,13,20,32,9,5,4,5,-15,-34,-14,-8,43,23,-26,-11,21),
	(-23,-24,8,-21,0,5,8,4,-24,-17,-44,-21,-11,-13,49,-21,5,-15,23,19,-6,29,47,-30,22,-7,-28,-12,6,24,-2,-4,33,0,-20,-17,36,17,34,5,-24,-21,6,-17,30,-11,14,20,18,25,-19,14,-4,27,21,4,47,30,29,7,33,-28,8,-4,-59,31,21,-6,16,-10,13,-5,42,15,-2,2,25,13,16,17,-9,31,41,0,-9,43,15,0,3,9,17,-2,5,2,11,7,2,21,9,-40,18,-16,-2,0,-4,7,-12,7,6,29,-15,-26,2,2,27,-2,1,3,1,15,-16,12,-14,17,34,-14,-20,17),
	(-40,11,0,-30,-5,-10,-3,31,-4,1,-3,-26,7,-40,56,-1,9,-13,-2,-8,-2,12,20,-19,6,12,-14,-9,-12,41,6,1,-6,-2,-25,-10,-3,-2,-2,34,0,-17,10,-18,9,-8,-3,33,27,8,-19,3,7,12,-1,27,24,17,-2,6,13,-23,-25,-7,-67,-2,-3,9,22,24,-17,-22,1,-16,13,37,0,1,23,18,-19,-7,63,38,-19,21,37,11,0,-2,32,7,-9,-1,-18,24,8,20,36,-16,2,-14,21,-35,-2,-5,4,-18,-12,29,0,23,23,-7,0,2,0,6,-20,-20,-6,1,-15,26,51,8,-11,-15),
	(-17,31,-9,-50,-2,-11,-12,43,-33,14,-13,0,3,-21,5,6,-11,-48,6,16,-1,20,39,-15,-15,14,-30,-38,11,-23,-16,-3,-3,-19,-33,-5,-1,-11,-10,7,-4,12,14,0,21,-5,-2,13,7,7,8,-14,-11,9,3,0,10,-5,13,-18,28,-3,-31,-9,-93,-18,-57,-3,27,-12,-1,-2,17,-12,25,11,23,-15,14,16,-36,2,23,46,20,-13,-16,25,7,-12,10,7,3,11,-7,-48,17,0,48,3,-4,9,-10,7,0,9,-16,-11,-13,-7,-10,22,11,12,3,-12,28,9,-18,9,-6,13,-27,21,28,-6,-29,-15),
	(7,8,-6,-53,11,-17,-13,26,-18,8,-27,16,-7,9,4,-16,-13,-11,11,-14,0,12,21,18,6,-19,-45,-40,-8,-7,8,-5,14,25,-13,-12,2,-5,-38,40,-18,9,11,-4,22,-11,10,10,32,-31,6,1,30,-9,8,0,2,8,7,-6,-18,-32,-36,-30,-52,7,-40,-4,0,9,-1,14,-13,13,1,35,15,-22,-12,-7,-16,-18,44,10,-18,-31,-12,-1,-4,13,6,-5,-23,-4,-15,-61,-12,20,40,-3,10,2,-30,-29,-18,-12,-12,-29,-45,30,-23,-18,12,-10,-27,-11,0,24,-48,6,27,11,-7,26,1,12,-9,2),
	(-13,28,3,-30,38,8,2,10,9,27,-1,19,-23,11,10,-10,15,9,-13,-6,6,-13,5,-19,-21,3,-13,-25,1,-29,-9,-5,0,-1,10,-7,4,18,-9,9,10,51,15,-14,15,-9,11,-7,27,-31,14,18,15,18,16,6,-35,-32,-13,-17,-26,-35,-20,-2,18,-1,-97,-1,18,3,5,-18,-64,16,26,50,2,-34,17,30,-2,-19,46,-33,-9,-31,19,49,-6,12,-20,-29,-16,13,-22,-50,10,5,13,-7,-6,0,-29,-7,30,-11,-27,-18,-9,15,13,-23,8,26,1,-27,12,11,-11,11,1,24,-28,27,32,12,-5,-15),
	(-6,60,-15,1,0,17,-10,-15,-6,11,-4,46,-22,-20,-4,10,9,-10,-18,18,-3,-10,4,0,-3,-5,-10,-5,-12,-22,-16,-5,8,-3,-19,5,-2,10,-38,0,21,8,16,-52,-12,14,11,1,30,-23,15,-24,21,-1,5,-10,-47,1,10,-13,-44,-45,6,-19,0,11,-73,13,52,-24,-19,-29,-79,8,18,32,10,-6,-21,11,-34,-41,14,-30,8,-5,-13,45,8,37,13,-3,7,20,-30,-33,-22,-8,-33,-33,21,-7,-33,-23,25,6,-3,-19,-27,0,14,-37,26,9,1,-14,1,3,-41,-4,1,8,-14,19,33,-8,-6,-33),
	(-29,18,13,-13,11,10,-23,-33,18,28,-1,64,-19,1,-13,13,9,6,-21,-13,15,-22,4,-4,-14,-17,15,-20,-8,-5,-16,-37,-34,-49,-9,-8,12,-14,-31,17,-6,3,-3,-41,9,9,11,32,-1,-2,33,-21,21,-16,24,-17,-35,5,-18,-2,-22,-44,16,-14,10,1,-8,-3,44,-24,0,-31,-61,13,-7,20,-10,-22,-13,17,-24,-43,16,-39,10,-22,-15,28,2,17,-1,41,-3,0,-20,-22,31,-11,-40,-4,-23,9,-7,8,6,7,-8,6,-14,-29,13,-44,29,27,8,-14,-6,-14,-16,8,-22,-21,12,-18,-4,-29,2,-25),
	(-42,30,-28,7,11,-14,24,-27,5,14,11,38,-15,-8,-20,-2,-9,20,-2,9,58,3,-13,-5,-2,-22,-13,-19,44,-16,-5,-24,-28,-17,1,6,-2,1,-33,17,-10,12,20,-8,-29,-25,18,26,-19,-9,20,0,4,-18,47,-11,-15,-1,18,19,-42,-29,17,-1,-10,14,-11,-32,20,-26,-10,-21,-32,21,11,18,-24,-39,10,25,-9,-38,0,-24,-6,-55,-5,20,-11,1,10,-9,24,5,15,-25,-3,-26,-38,-42,1,5,-49,19,40,13,-28,1,-13,-19,-20,-15,-1,-3,-37,-11,-4,26,-39,-26,0,2,25,21,19,3,-18,-41),
	(5,-24,-26,20,-16,40,37,-17,16,3,52,-22,19,-16,-7,35,24,-3,-1,0,31,-41,16,-9,-35,29,-33,12,31,-43,29,-21,18,-38,34,-61,47,-21,-15,-14,-42,-2,93,60,-37,-65,26,52,-70,-23,-21,-21,-25,-11,62,9,-10,30,-25,17,-56,22,36,-2,14,-16,25,-14,1,-10,-13,-14,9,36,-19,0,42,0,44,11,-12,-19,34,2,-21,-58,38,-14,-9,-23,-31,-75,0,31,-28,2,-1,36,-57,18,30,10,-41,-27,22,38,-47,7,-16,-10,-50,24,-2,-66,-51,4,13,63,-10,-14,72,56,61,0,54,-15,14,-44),
	(29,-57,-39,-5,43,-12,9,33,22,-26,41,-32,35,13,-21,7,15,14,-21,12,22,2,15,-2,-37,-11,-14,24,21,7,22,-27,-9,-23,64,1,16,5,1,20,-14,1,15,28,-31,2,3,-2,-24,-18,-9,9,-34,14,29,35,8,28,3,-16,-13,18,5,-3,26,-17,11,-31,5,-20,-13,1,24,17,-14,-12,10,4,4,22,-33,-26,9,6,-12,-32,5,-7,-40,-5,-52,-65,-48,10,-9,-27,11,-4,0,20,10,-34,-42,-22,11,-12,13,17,-23,5,-1,28,-32,0,-19,7,-52,50,16,12,14,23,4,3,4,-32,21,-4),
	(0,-62,-20,16,-39,0,37,10,12,9,38,-15,29,-3,-26,21,12,61,-59,28,25,2,-13,3,21,18,-15,8,-16,-10,38,-40,30,-28,22,-5,9,42,-27,-36,-18,-15,37,42,10,-34,29,-24,-48,-32,31,55,19,5,26,-34,-34,2,-10,-9,22,18,55,-27,-14,0,35,6,15,-27,12,40,24,35,-27,-31,5,9,-50,-10,-31,28,35,-24,13,-19,-16,-30,-30,-41,-54,-9,-13,27,-1,-24,24,-3,-41,-7,26,-28,19,21,-2,34,-47,-22,-25,20,-40,29,-12,-28,5,9,20,28,-5,21,21,42,61,14,16,-7,17,-28),
	(-1,7,-11,11,-9,-27,0,0,22,2,9,-13,15,22,40,11,-39,-20,-16,31,36,14,-17,1,24,-25,-14,5,14,-3,-8,4,-20,-7,30,-36,25,-14,-27,29,-4,3,6,27,-2,-9,-19,-13,11,21,8,-27,13,-10,32,14,-9,19,8,-11,12,-12,36,0,-1,21,-11,5,13,1,1,-19,44,41,32,-6,-26,23,19,-6,-8,-19,0,-14,-8,-14,5,-26,-8,9,-32,-4,31,-1,32,-1,-15,14,-31,23,-11,-28,-27,-24,0,-43,7,-3,-34,-18,7,0,-20,-11,-6,13,21,30,-2,3,-18,13,17,29,0,-8,6,-7),
	(5,-16,2,11,9,-11,4,17,-1,-4,14,12,-18,11,-22,-17,-4,-2,2,5,-11,11,28,-9,-10,16,-4,10,32,0,0,27,-13,5,-20,19,-20,0,5,-3,17,3,1,4,-5,28,-10,-30,8,-9,16,2,-26,13,33,-16,7,10,7,5,-10,31,16,-14,6,-19,-11,-8,-1,-3,-2,-5,-10,34,3,25,-34,29,-29,-3,2,9,6,1,33,-17,-4,1,1,4,-14,-3,-22,-7,-21,17,1,0,-10,28,-31,-16,30,9,-11,-19,16,6,20,-14,0,-9,22,17,30,29,6,-8,3,4,-5,-32,-4,-19,-11,-11,-23,11),
	(4,0,31,-28,23,-1,-27,3,39,33,-35,4,-4,-3,25,-4,25,5,15,12,-32,10,33,-45,-24,-19,-4,-17,61,22,-37,15,-11,-24,-3,18,1,22,6,0,0,-10,-1,12,13,-11,24,-15,0,28,17,29,-27,-19,11,26,14,-6,-24,8,-16,-17,-23,24,-22,-37,-21,-23,-8,2,-5,8,-31,-1,18,35,-27,-7,18,21,-9,-10,-6,25,17,28,16,19,-8,30,15,-8,18,-15,-18,-7,-22,1,5,3,5,-46,-18,-5,3,-18,13,7,28,7,-2,-33,23,0,17,-8,-13,27,-24,36,-28,0,-8,24,25,-35,-45,23),
	(18,0,-33,18,8,18,-41,16,40,-16,-58,-12,-14,-44,-28,-24,31,-6,19,38,-19,-51,4,-46,-36,48,-5,21,18,3,23,37,27,-7,-22,-12,-31,74,-15,40,38,29,-19,-39,61,23,34,-2,1,1,15,38,-64,29,41,12,-19,0,-40,1,16,44,14,-34,8,-31,-59,-2,-30,-38,38,36,-40,-26,52,20,-25,20,-14,28,-24,26,38,-21,11,-33,-7,54,-5,-4,13,-10,-27,-12,-66,-15,2,56,24,0,2,-3,-12,-11,-37,-6,-53,-30,-18,-35,-25,1,43,39,24,16,38,29,0,45,16,-43,-16,-37,15,-41,-22,1),
	(5,-10,-46,8,7,4,-24,5,2,-10,-71,-39,-19,-57,-5,15,13,6,3,30,-28,13,-10,-32,-2,-13,-2,-2,10,18,10,-13,22,4,-11,-18,-4,56,-48,42,19,13,0,-17,10,7,39,10,-10,0,-12,46,-10,1,18,19,-16,-15,-5,-1,2,-7,27,-37,-11,0,3,-1,-41,25,-18,-3,-14,-45,15,-43,11,-3,-5,31,-21,24,28,-21,0,-11,10,20,-5,9,6,-27,-14,-32,-32,-1,21,26,34,-34,22,-45,-4,2,10,-11,-26,-26,-45,15,-17,-17,-13,20,20,-27,-16,14,-18,29,13,3,-7,-43,30,-21,13,-15),
	(0,-7,-10,-1,18,0,0,-5,22,-2,-78,-37,-14,-31,-8,2,-12,11,-15,-2,-11,19,-16,-40,-11,0,-27,31,3,-21,30,-11,33,6,-26,-17,10,17,-32,11,-2,-10,3,-48,38,-7,-20,19,3,2,19,45,-16,-11,14,7,-14,16,-15,0,11,12,-11,-8,-13,-8,13,-18,-19,10,0,9,28,-15,2,-26,36,16,-5,5,-21,40,25,-33,-14,-2,-68,27,-24,-51,-21,-18,-3,-20,-38,-14,-6,1,43,9,-2,-19,14,13,-33,17,-45,-17,-45,17,1,-35,14,18,35,-32,-20,-13,-26,-16,-28,0,-24,-32,-1,-14,16,-1),
	(18,8,-34,-28,-12,24,-1,-39,-5,-33,-51,-19,23,-48,3,12,-8,24,-14,-9,8,-2,9,-11,17,1,-34,11,-3,-14,22,-9,18,-21,-17,-16,-2,37,-49,0,0,-10,-18,-72,47,2,-25,40,30,-25,20,30,0,-12,23,4,-15,8,-14,0,-4,6,-7,-31,-28,3,23,-27,-29,-24,10,-31,21,-18,2,-31,34,-6,-15,-6,1,64,7,-55,-4,-38,-110,4,-21,-34,0,7,4,1,-48,-19,-2,16,60,-15,8,4,-5,-16,-8,4,-10,-21,-67,-6,9,-30,5,-2,0,11,6,-6,-47,-36,8,6,-27,-77,-5,-7,-17,-15),
	(9,42,6,-4,-11,13,13,-60,-8,-6,-17,-57,30,-4,12,10,-10,24,-21,-6,-7,-1,31,10,6,0,-38,-2,27,-10,42,-28,28,-5,-28,-7,34,19,-50,0,-17,-22,-52,-69,2,-15,-31,15,8,-9,8,6,-2,-24,1,4,-10,12,-17,-7,25,24,5,2,-32,0,43,11,-3,-6,-10,-9,33,-19,-5,-17,42,-7,-6,17,-17,35,42,-8,-10,-26,-72,0,-23,-32,16,9,-19,-13,-20,-56,-4,33,26,12,17,-65,-5,8,-1,3,-6,-37,-91,27,7,2,15,6,-18,16,0,-22,-44,-12,6,28,-41,-86,-3,10,20,-15),
	(27,51,-12,3,-17,-10,32,-27,0,16,-9,-41,26,29,-19,21,30,12,-11,16,-11,24,26,-10,-3,23,-19,-17,-9,-31,25,-21,6,1,-3,-23,-6,8,-57,-8,-55,-9,-61,-39,9,-17,-9,-5,4,3,18,-10,13,-36,13,-22,0,-13,27,3,14,28,9,-7,-17,26,0,-10,-25,3,19,7,38,9,-26,-40,0,-1,13,20,-12,-12,22,-2,-23,4,-112,-29,-11,-32,26,5,-3,5,-43,-46,15,8,30,-16,-1,-36,-5,10,13,18,-8,-36,-66,-2,12,-8,-9,8,-33,30,0,-23,-50,-51,-6,25,-46,-74,6,-8,1,-31),
	(34,40,-16,-2,-9,24,13,-18,20,6,6,-38,16,29,-40,2,3,6,9,2,7,19,0,41,1,29,-16,-2,-12,-49,17,-10,-13,-16,8,-4,-20,15,-10,-25,-39,-6,-38,10,-4,-15,25,-34,0,-8,43,-6,20,-27,-22,-17,-31,-16,21,-18,-3,18,7,22,-22,13,-2,3,-2,-4,7,-13,16,-19,-15,-44,15,-8,0,-4,-3,-28,11,17,-23,-7,-96,-25,9,-19,-15,-21,-18,21,-9,-50,-8,-15,6,-18,34,-6,15,1,19,7,-27,-23,-48,5,8,-8,0,2,-8,37,-8,-48,-42,-62,7,27,-28,-134,0,-14,23,-3),
	(38,50,-12,0,-10,-2,15,-20,15,-8,34,-16,11,44,-64,-3,9,17,42,5,13,-27,26,0,-17,6,38,16,-37,-35,28,-12,0,-28,5,-54,-10,-14,-21,13,-46,-1,26,45,25,-33,64,-41,-9,-3,6,-14,22,-14,-13,7,-26,-7,5,-12,-9,25,7,13,-51,9,27,22,-5,-29,22,12,28,15,-43,-43,32,-4,-22,2,-12,22,8,-2,-16,-5,-109,-30,11,-14,-22,-3,15,3,19,-26,-8,-11,-12,-24,10,1,15,0,11,33,-30,-4,-32,-17,-20,-8,4,-31,19,8,4,-43,-38,-34,0,17,-18,-109,21,3,14,-19),
	(26,10,-29,11,17,-2,-31,20,-23,1,43,1,28,52,-41,4,-2,0,19,3,16,-48,10,20,3,8,18,17,-8,-26,5,8,-6,-4,9,-32,6,9,15,-5,-41,17,33,20,13,-43,42,-62,4,-25,-10,0,-4,-42,-24,-10,0,18,19,-16,-26,14,1,13,-20,8,1,11,-3,-7,15,-11,-1,-19,-28,-47,33,-4,-35,19,-5,19,-20,1,-29,9,-70,-26,17,-16,-42,-26,9,-21,43,-17,-24,23,8,4,10,-2,-40,0,11,21,-16,48,-42,-17,-2,-8,0,-19,18,16,22,-35,-13,-36,-21,27,26,-100,2,1,-13,3),
	(23,14,-31,-13,-10,-3,-11,-7,2,-17,54,7,9,24,-43,4,-9,-21,47,2,-18,-40,14,0,-22,13,40,-3,11,-12,11,2,-14,-27,42,-31,-6,15,23,-14,-70,22,62,0,43,10,35,4,-9,-13,-47,-5,-32,-69,-30,0,2,4,-21,-11,-20,4,0,27,-15,1,0,1,2,-21,21,-12,13,-33,-52,-57,19,3,0,9,5,18,14,36,-29,-11,-134,-2,50,-4,-54,-43,-3,19,13,-40,-31,18,32,24,2,39,-11,-1,0,5,-11,29,-21,-38,-25,-15,38,-20,1,-26,24,-40,-26,-36,13,16,39,-15,-3,21,9,-14),
	(34,-7,-17,10,19,33,5,11,-17,-24,33,1,18,53,-25,-4,17,-3,13,-12,-12,-68,-21,15,-23,27,-4,11,31,-31,10,-3,-21,-17,19,-24,-11,20,22,-13,-80,38,11,14,17,8,31,8,-7,-11,-57,12,-7,-49,-12,24,12,-8,10,-6,-21,0,-8,0,-12,-17,3,13,5,4,11,10,10,-16,-5,-34,22,-6,9,8,12,0,11,2,-23,-3,-133,7,36,-1,-18,-38,17,23,21,-45,-29,4,41,0,11,44,-23,-24,19,14,5,21,0,-17,19,-26,4,2,15,-2,-3,-23,2,-41,1,-15,31,46,21,-21,-25,18),
	(0,-6,3,-20,-18,31,4,0,-6,-35,11,-25,31,14,13,-2,26,-12,-10,15,-11,-51,3,-38,-5,19,-28,-17,7,-31,25,10,-32,9,12,-36,24,-4,11,10,4,-5,2,3,-2,35,18,27,10,2,-17,-5,-15,-10,-6,5,34,-14,7,7,-7,0,2,-12,12,0,26,1,-32,19,2,-21,50,-15,-11,-16,18,12,8,2,-3,3,26,9,-21,16,-61,-15,-19,-22,32,-56,14,-9,-18,-15,-46,2,1,0,-5,10,-26,-25,-32,-13,11,-7,-7,12,9,-37,-5,-19,1,-10,1,-6,24,-23,-12,-10,2,70,24,-32,-19,0),
	(14,-35,18,7,-17,-8,0,-17,-15,-1,1,-51,12,-33,44,1,3,-1,19,20,-8,-58,9,-11,22,11,-34,-13,21,-20,5,15,4,12,5,-28,25,32,-2,31,22,-7,1,-28,21,5,12,32,9,9,-14,12,-29,31,25,12,24,14,10,-13,4,-10,-17,-13,-8,-2,16,10,-36,-18,17,11,49,7,15,18,-19,8,0,11,-7,-28,62,-5,-2,19,-22,-1,0,5,47,-18,-33,-11,11,10,-22,-11,16,-8,11,16,6,1,-46,-2,4,18,10,17,-16,-21,-5,19,-2,4,-15,2,-6,-2,-27,-4,2,54,49,-22,-6,25),
	(-5,-25,18,5,-16,20,-12,-15,-18,10,9,-53,12,-24,35,15,39,-8,-1,8,-15,-24,35,-37,-5,10,-3,15,10,25,2,7,22,3,-19,-12,-3,21,0,29,19,-23,-2,-14,26,-21,22,4,-1,16,-18,5,-13,2,-6,-17,12,-8,0,10,13,3,-13,-2,-45,0,44,16,4,-16,-17,13,29,-18,-13,35,13,11,-9,13,-11,18,38,-33,-12,26,34,-4,-10,-10,12,-2,-2,-37,16,9,-1,-16,-6,-15,1,10,32,-2,-9,-1,13,22,22,34,8,-10,28,11,12,-9,11,6,18,4,-2,13,-21,44,61,-11,9,4),
	(-22,11,-13,-6,-15,10,8,-5,-9,-1,-10,-17,16,-26,29,1,9,9,31,1,1,7,9,-26,2,-2,-7,-3,-3,11,10,23,32,17,-24,-13,19,20,-5,-3,28,-24,26,-9,3,-23,18,44,-5,-4,-36,-9,-11,30,-7,-22,23,14,-3,13,8,-28,10,-23,-83,13,3,3,17,-17,0,0,36,13,21,37,-6,-23,5,-2,17,-4,29,2,-1,7,37,10,6,19,19,21,-8,-15,4,23,5,11,8,-26,0,-27,40,-11,-24,-24,-27,21,-10,4,-22,14,3,-8,-7,1,25,-4,0,11,-26,13,-41,27,42,-17,-5,13),
	(-18,19,-24,-12,-14,-10,7,15,-4,21,-10,-7,-12,-42,3,0,10,-5,-9,-2,-4,22,49,-2,-12,21,2,-7,19,43,-17,11,22,5,-23,-2,15,-2,10,6,-8,-11,25,-14,7,-29,45,15,7,15,-35,-8,-4,0,9,-22,16,-9,4,-11,-3,-26,25,-3,-78,-8,-16,-11,10,12,9,-15,26,1,16,7,16,-31,4,6,11,31,46,-5,-9,3,3,8,12,2,15,20,-21,23,12,20,-5,22,23,1,-2,-5,9,-13,7,-15,-8,-13,-12,7,-11,22,-8,-4,-8,7,-14,7,-20,10,2,-3,-16,35,35,-9,-7,-2),
	(-15,47,-20,-13,-30,-1,-26,53,0,13,-4,16,-12,-22,-2,-3,-14,-18,3,18,-4,-14,2,-26,9,-3,-8,2,19,-6,-3,-9,16,11,-24,11,1,26,11,36,16,-24,13,-27,24,-32,4,5,29,-22,-53,6,-29,37,0,-5,9,-12,12,-18,29,-4,31,-7,-55,4,-74,-6,20,-16,-1,14,-1,-5,19,39,-15,4,10,-22,-31,39,10,8,-11,0,5,15,-8,21,-7,39,-5,2,-23,-21,-6,-7,24,-17,-11,-24,-2,-6,-13,-22,-1,-20,-25,17,-7,-7,15,-10,-18,-16,19,-22,-16,26,-14,6,-38,23,24,7,-31,1),
	(-10,24,-20,-37,4,18,-18,20,4,-3,-12,26,-8,1,4,-6,-13,-14,-13,16,0,-7,-8,-21,6,-4,-44,-17,-6,-41,-7,-16,2,25,-9,6,8,3,-9,14,20,6,1,-28,-13,-5,-4,5,17,9,-3,14,-4,15,3,2,-17,-15,16,-17,-5,-1,9,-14,-59,11,-74,-6,25,25,-14,3,-41,29,24,31,19,-12,-11,0,-10,17,24,-28,11,-19,8,24,8,21,-3,-14,-6,24,-21,-66,-7,-5,-14,0,18,7,-42,15,0,-7,5,-27,-40,-13,19,4,23,-11,0,-7,-21,-2,-55,0,-2,5,5,9,-7,-1,4,6),
	(13,31,-22,-6,25,11,-17,33,-32,2,-5,14,-32,-21,-11,-11,4,3,-12,-2,6,-19,22,-20,-4,-20,-17,-13,26,-13,10,-13,-22,3,11,-13,5,3,-17,18,30,31,-10,-24,13,20,-10,16,0,-18,22,1,5,19,7,12,-33,1,0,-7,-16,-15,31,-14,-16,-18,-85,-6,21,-19,-10,-3,-90,28,6,35,4,-27,-21,17,-9,5,20,-62,-12,-6,-7,26,22,13,-10,-17,-7,14,-11,-70,-5,18,-12,-2,-5,-36,-32,-21,2,14,-1,-25,-23,0,-3,-28,1,23,-10,-27,-14,33,-17,31,20,11,4,-10,12,-11,9,-2),
	(0,42,-17,3,-13,4,-1,-4,-16,27,0,39,-1,-25,-19,17,0,-5,-5,28,15,-13,24,-32,-22,-19,-22,-25,-10,-31,-10,-28,14,-45,-8,-6,14,26,-25,-7,8,-7,-9,-42,-20,-15,2,6,-14,0,30,-14,11,3,26,-21,-63,-3,15,17,-24,-7,34,-5,0,4,-65,-5,2,1,24,-15,-56,12,13,29,-20,-33,-13,-10,-33,-27,12,-75,17,-11,8,38,3,15,-16,9,10,16,-3,-20,2,-21,-29,-12,15,-27,-15,15,-10,8,2,-12,-34,-39,-3,-13,-12,6,10,7,-4,0,-49,12,-4,0,15,-3,18,-8,-6,-10),
	(9,4,10,-19,-31,26,7,-29,11,-8,12,40,-21,-7,-34,-5,12,-7,-7,-4,21,-28,11,-6,0,20,21,16,-1,-29,17,-33,4,-53,2,10,-13,22,-46,-8,13,5,13,-5,-9,-22,22,31,-19,-15,49,-9,-4,-14,18,-35,-32,2,-31,0,-42,-11,28,1,22,-31,-39,-4,4,-16,-5,3,-19,-24,3,9,15,-34,-25,2,-33,-7,21,-67,2,-59,-19,26,25,-20,18,-7,-3,-16,-23,-50,16,5,-38,-31,-11,-8,-21,3,-22,33,-18,-12,-30,-7,-19,-29,16,28,-24,26,-24,5,-46,1,8,0,23,-20,19,0,-14,-24),
	(-2,-2,-20,-9,-7,3,15,-25,10,-7,27,18,24,-14,-21,25,-16,18,-32,-15,0,-37,-2,-2,-16,-1,28,12,4,-42,3,-15,-13,-40,34,-21,10,25,-26,-8,6,-15,12,5,-3,-42,-32,37,-1,-22,6,3,0,3,38,-24,-24,-3,-37,-9,-37,13,15,-24,-1,-31,-9,-35,-20,-18,-17,-13,-31,-23,0,-1,17,-17,-27,-18,-8,-6,15,-70,13,-46,13,7,-33,-38,34,-18,0,23,1,-51,1,-35,-46,-19,19,17,-74,-20,-2,0,-34,-31,-33,-28,-2,-23,-22,-12,-44,13,-24,15,-32,-24,12,20,27,-5,45,-1,15,-58),
	(29,-19,-14,10,3,55,0,-2,42,-23,2,-41,13,-7,-3,36,17,27,-47,4,29,-23,-1,-13,-36,49,1,12,30,-11,14,-5,-15,-43,49,-52,5,9,-27,-34,-16,-21,48,57,-47,-52,9,30,-49,-29,-5,-38,-29,21,42,-12,-24,-3,-31,1,-28,9,29,-16,23,-57,0,9,34,13,38,-15,25,3,2,0,12,28,-15,-8,0,1,47,-39,-2,-26,19,6,-23,-13,-7,-56,-11,44,-9,12,-17,9,9,27,33,-31,-38,-43,12,7,-45,6,-41,-23,-18,20,-18,-49,-33,51,3,37,5,-1,27,37,17,-13,59,5,26,-15),
	(1,-56,-12,7,16,9,-12,4,31,-20,4,-25,45,13,-12,11,-1,30,20,17,13,-5,-28,23,-37,4,-4,5,49,13,26,10,4,-5,42,-6,30,-20,-3,35,-40,13,39,-9,-43,-2,16,11,4,-9,-25,-12,-20,13,37,14,2,26,12,-13,-23,36,32,-4,38,-15,16,-41,66,-22,-5,4,4,57,-26,-22,6,-27,15,21,-13,-22,-4,38,-17,-6,-12,-12,-25,0,-23,-7,-2,8,22,-12,-23,-1,-11,10,-12,-47,-19,-34,29,-16,20,2,11,-16,31,28,-40,-10,24,3,-9,34,37,-14,37,-11,2,32,8,-55,17,7),
	(51,-53,2,6,26,27,41,56,32,-18,24,-33,45,2,-9,20,45,25,-17,24,19,14,-10,-21,-37,51,-6,28,28,-21,28,4,29,-49,33,15,19,35,5,0,-45,-8,48,23,29,-3,-6,1,-28,-7,-18,42,-32,33,47,-13,-9,-10,-18,6,-8,31,25,25,34,-23,0,-10,3,-14,26,24,34,26,-29,20,43,-9,3,36,15,6,46,23,-10,28,8,36,-12,-2,-11,-16,-27,-3,-9,-13,-6,8,-25,-21,48,-9,0,-28,8,33,-32,0,36,-7,-30,31,16,-13,-19,18,12,39,-5,36,29,27,23,-13,62,-24,44,18),
	(6,0,-11,-14,-1,3,-19,-4,-10,14,2,-20,-8,-13,-18,-18,-16,8,0,-17,18,-8,0,17,12,5,17,3,0,7,-5,-3,4,-4,2,16,0,22,7,14,11,18,-15,-3,9,-12,-7,4,-1,-7,3,13,15,15,-17,9,-7,-11,8,-16,6,13,8,21,-12,16,-15,-16,0,-11,-9,-7,21,-17,3,-18,3,0,16,-1,20,-15,14,23,16,16,-6,-7,9,20,-16,-10,0,16,-9,-16,-15,-1,-6,0,-16,-2,-13,-5,-18,-17,-16,-21,13,-7,1,-9,-15,5,0,2,-12,-9,-12,2,18,-7,-13,-15,2,15,9,6),
	(-35,-2,0,18,-4,-28,18,14,20,23,14,-17,19,7,31,9,-16,10,-4,10,34,-4,-6,7,9,-13,-21,17,-8,3,-2,38,16,14,9,-7,37,-34,-28,16,13,16,18,6,-13,17,17,-8,4,32,46,-14,18,18,16,0,-19,18,18,9,50,27,0,-26,-30,1,35,-10,-5,19,-8,4,11,21,-3,-3,-22,-11,15,-1,-14,-24,0,1,-15,17,21,-6,-15,23,3,-23,20,21,37,0,-9,11,12,21,-18,-31,-12,-41,30,-9,-37,9,-33,-13,13,6,-39,-2,-1,7,0,17,-12,26,1,15,19,49,15,0,-7,-23),
	(-17,19,6,-9,3,-21,-27,9,-23,3,-12,20,-26,36,0,-10,0,15,12,1,10,38,-16,-16,-11,-22,-36,-7,0,-6,21,-15,-5,23,18,-11,14,-5,19,3,40,18,-32,-13,12,-16,0,-6,8,0,-1,-14,3,5,2,-9,28,7,-30,-19,-9,-2,-29,-29,-45,6,-5,1,6,-9,-42,-18,-18,-21,-3,-10,6,-1,-6,-4,7,-6,-16,-8,-28,-6,43,5,10,-9,18,-8,14,-21,-26,-16,-12,10,0,4,-9,-55,-22,-42,10,-26,-8,-3,-1,0,15,27,-34,-20,-1,-34,-21,25,-12,-12,10,5,-2,22,11,24,-12,10),
	(-6,36,-13,-21,24,-8,-48,2,17,-21,-11,-10,-16,-30,-48,-30,48,-11,5,4,-27,-63,14,-44,-10,1,-12,14,5,-7,-5,-4,33,24,-8,16,-7,23,-5,32,18,-7,-12,-24,40,24,-14,2,10,22,-21,65,-47,-9,13,28,8,-20,-14,19,-6,26,19,-17,5,-39,-71,7,-51,-4,2,6,-43,-26,10,27,0,13,-11,39,12,28,43,15,-2,14,17,35,24,-8,16,18,-12,-33,-52,12,9,0,47,7,15,-37,-12,-38,0,-8,-27,-48,-5,-18,-28,-6,30,25,0,1,-18,44,-13,39,12,0,-4,-63,37,1,-10,12),
	(-8,4,-62,-4,-16,13,-26,4,0,8,-22,-9,7,-32,-12,-12,41,1,23,-5,-4,24,-14,-47,0,8,-8,-9,21,4,25,4,27,5,-24,-27,20,46,-10,19,3,12,0,-29,30,-21,-6,18,18,-6,-1,20,4,17,9,11,0,-5,9,-4,-17,0,17,14,8,-5,-1,-4,-20,23,-11,9,9,-8,11,-8,16,16,10,11,-10,47,46,28,-21,-4,0,31,-26,-18,38,12,-12,-5,-56,38,8,-2,17,0,10,-55,-13,-3,-3,10,-41,-22,-28,0,-13,-15,-11,25,6,-18,-21,25,-8,-12,10,10,-6,-24,24,-5,17,-8),
	(-14,3,-40,0,18,2,-23,-14,27,-35,-23,1,-5,-56,-23,-18,17,-7,-8,26,-9,29,4,-29,13,16,-16,4,7,18,7,-5,20,9,-21,-13,19,19,-28,27,17,-4,0,-60,34,-24,-7,31,12,5,7,29,8,-5,12,-9,-8,23,-18,4,0,1,-22,-20,-7,3,21,-29,-37,3,-1,10,41,-35,29,-11,-7,22,-29,26,-18,45,36,13,-3,-25,-51,19,-29,-24,2,24,-6,-7,-36,14,2,14,24,13,22,-8,1,17,-41,16,-11,-35,9,16,-1,-29,4,13,6,0,-8,2,29,11,0,0,-34,-83,-5,-25,-3,0),
	(-17,6,-51,-11,7,6,0,-51,23,-1,-13,-21,21,-39,11,-9,6,-3,-7,16,7,19,6,-20,21,16,-54,12,-7,10,34,9,-13,-13,-38,10,-6,3,-14,25,7,13,-37,-57,33,-14,-54,25,24,-2,20,25,14,0,25,-5,-15,-10,17,-10,2,17,-11,7,-24,-10,-2,-26,-57,3,-17,-9,38,-36,38,-25,22,6,-20,5,-19,18,12,-5,5,-20,-39,5,-10,-42,4,0,-27,-6,-53,5,-10,6,32,7,11,-14,3,18,1,19,-35,-11,-40,3,-5,-1,-4,26,-2,-13,2,-12,-21,-10,-5,11,-21,-88,-36,-7,5,-17),
	(-4,19,-53,19,0,3,30,-52,0,-25,19,-6,13,-24,-15,6,21,20,19,27,-18,18,17,6,-23,21,-36,-3,20,-13,-3,-11,6,-20,-20,-23,-6,8,-26,-11,-23,-5,-41,-54,16,-2,-13,-35,-27,-7,37,3,-2,-34,11,2,-4,3,4,-3,16,32,3,1,-38,-4,18,10,-81,8,-4,22,26,-27,0,-33,-1,7,17,-2,-26,0,26,13,7,-37,-70,8,-9,-25,15,5,-10,6,-44,-38,-14,-11,60,2,22,-45,5,-24,23,20,-43,-19,-54,27,-7,1,-5,-7,-26,27,-8,-12,-35,6,10,-10,-37,-64,-22,-8,3,-13),
	(-3,20,-39,16,-23,-11,42,-31,13,0,21,-26,22,-49,-19,-13,-4,-1,23,7,6,28,31,19,13,15,0,-4,0,-20,21,-5,1,-23,24,-19,4,-2,-47,10,-19,-4,-84,-41,18,-9,15,-14,0,0,48,28,33,-8,27,6,12,22,0,-3,22,17,33,26,-61,0,5,16,-60,6,-18,14,18,-39,-16,-20,2,2,1,22,12,4,14,-25,-3,-26,-81,-8,-19,-29,8,-7,-13,-10,-43,-51,-16,-7,44,6,8,-10,17,-13,25,6,-32,-26,-75,1,-5,5,4,-20,-4,25,-19,-3,-43,-1,29,1,-41,-59,9,11,-10,-8),
	(-23,50,-69,18,-12,-11,19,-11,3,3,28,-10,19,-4,-47,-5,11,3,22,1,2,-18,13,21,-5,-5,28,6,0,-24,4,6,-9,-4,31,0,-20,0,-22,11,-16,11,-38,21,-4,-26,49,-4,-21,7,7,-10,27,-32,5,-17,-20,-1,-6,11,-9,23,34,16,-42,2,10,-1,-57,-8,19,31,35,-40,21,-30,24,6,-1,0,12,-28,9,-12,-5,-26,-80,15,-4,10,-2,-6,-25,33,-12,-72,-1,-7,17,22,-16,-31,-9,6,10,2,-48,-11,-78,0,-18,0,21,-8,-20,8,21,-25,-52,-10,-10,32,-9,-103,-6,3,22,-28),
	(-1,47,-62,18,-8,-5,9,0,8,-7,35,-7,28,-1,-65,11,19,-13,38,-7,3,-48,38,26,7,18,23,13,-35,-37,13,-1,23,0,20,-22,-25,-12,-18,-16,-47,-3,22,49,15,-40,32,-23,-15,-19,-27,12,15,-50,30,-14,-11,3,-4,14,12,16,-3,10,-29,13,22,21,-53,-37,10,0,34,0,-8,-1,27,11,-31,10,2,6,13,-29,-17,-10,-81,7,5,-1,-32,-28,7,37,9,-29,-9,7,25,9,13,-17,1,-7,34,13,-28,28,-79,-38,-6,23,22,-13,-33,11,26,-24,-52,-21,15,27,4,-72,9,2,21,-9),
	(-9,31,-64,-11,0,3,-32,7,-28,9,50,-32,2,9,-67,-6,6,-31,32,-8,-24,-38,21,8,-28,10,18,22,-37,-18,-4,-21,2,-13,47,-48,-1,-12,-20,-11,-40,17,23,30,22,-39,27,-25,-10,-15,-30,-11,0,-42,11,-29,-6,4,-4,-9,-9,24,21,-11,-31,-10,-3,-6,-60,-33,-11,-6,14,-44,-33,-5,28,7,-22,-13,-7,9,9,-15,-41,-28,-51,20,27,-20,-34,-41,3,14,28,-66,13,-9,11,-3,6,14,-30,-37,9,20,-23,49,-36,-45,-33,7,-10,8,-46,28,-8,-26,-23,-20,3,17,63,-34,17,22,3,-13),
	(7,0,-39,8,-15,-8,5,36,-45,-1,41,-5,16,37,-20,-6,0,-1,5,16,-7,-44,13,11,0,2,13,-7,-13,12,-7,3,9,10,12,-56,7,-22,-30,-7,-33,-8,54,20,-10,-23,30,-8,10,-21,-29,-9,-9,-47,18,-10,-6,9,-4,-2,0,47,5,0,-15,11,8,2,-45,0,3,-1,61,-23,-25,10,21,-3,-3,24,-10,4,-15,7,-2,-29,-92,35,7,-1,-30,-25,19,20,16,-54,12,-10,41,18,-18,34,-26,-26,1,-14,-25,43,-62,-29,-24,-1,14,-14,-46,24,22,-2,-32,0,10,0,74,4,-3,20,-10,-17),
	(-6,-13,-15,2,11,23,13,13,-1,-8,42,-12,0,26,-5,21,-5,-27,16,17,4,-47,-18,-6,-11,9,-3,-11,-11,27,-5,19,12,4,32,-49,-2,15,-32,14,-24,-4,33,28,-3,26,-8,32,0,-30,-2,-10,-33,-8,15,-8,-15,-7,-4,6,-10,45,10,-3,13,-20,0,12,-58,6,-6,-2,40,9,-18,3,5,10,19,19,-16,-7,-14,7,11,1,-97,3,-4,-4,-19,-32,-8,3,9,-31,4,-8,34,4,-13,59,-25,-8,-10,23,-17,22,-47,-21,-23,7,1,2,1,16,4,28,-17,5,-2,-10,23,38,5,-7,-8,4),
	(-9,-40,1,6,-10,2,-1,-27,-31,-13,35,-31,1,-37,56,0,17,-28,-11,14,-1,-48,-30,-15,18,-13,-34,9,21,0,10,8,-26,17,-15,-9,22,10,20,2,16,-2,15,5,-1,36,18,15,-7,17,-10,8,-37,15,25,10,-4,0,9,-12,0,12,-2,-18,23,1,34,2,-38,15,1,11,23,12,16,28,15,-5,5,20,3,-29,38,-18,2,2,-40,17,12,-7,40,-43,7,8,-20,7,-22,-14,15,2,22,5,-7,-19,-38,-24,1,-3,-30,2,0,-8,-11,-14,-18,9,19,2,0,-1,-4,-36,10,41,27,-31,-15,-7),
	(-14,-43,23,-12,5,34,11,-2,-23,-36,30,-20,27,-70,36,-8,27,6,19,13,-3,-41,11,-20,-23,-8,-23,0,10,11,5,11,-16,2,-7,1,21,10,12,7,32,-22,19,-3,13,11,26,5,-7,-13,1,-20,-48,7,24,12,9,-2,-18,3,7,1,16,-13,-36,-11,36,23,-17,-11,-6,4,40,-22,21,35,-13,-15,-5,15,23,-28,24,-41,14,30,-7,10,6,1,61,-17,-21,-24,9,-4,20,-29,39,-9,36,-4,15,12,-21,-9,6,4,9,13,-1,-2,-1,16,4,17,-11,9,12,2,9,7,-7,55,19,-27,0,8),
	(-2,-23,17,5,12,-1,-6,-62,6,-9,0,-16,24,-53,11,0,20,20,2,11,-8,-23,27,8,-3,22,-4,3,28,4,-10,7,15,-9,-12,29,-11,11,18,2,43,-24,5,-4,18,-15,-1,24,2,9,-10,0,-32,16,-18,-4,13,0,-5,-12,22,-22,16,-7,-49,-11,35,24,-12,-20,-1,20,-10,10,7,19,-1,14,-6,-22,10,16,41,-29,11,-6,34,5,4,-1,31,-16,1,-1,-17,9,17,-35,43,-18,27,11,32,16,-14,-16,-12,11,6,9,-21,14,5,0,-6,16,16,15,10,9,-4,10,-43,30,9,0,1,33),
	(-11,4,-19,-3,-6,7,-24,-19,10,30,14,2,-16,-21,3,22,-4,28,18,22,-21,30,25,-15,8,9,-7,-14,-6,4,24,20,9,4,-29,-6,8,9,-11,25,27,1,-3,2,0,-18,23,41,1,14,-31,16,-5,9,-16,-8,37,6,0,-5,3,7,3,-7,-60,-2,-12,23,-9,-25,26,10,-8,-5,2,-12,0,0,-1,-15,1,-1,30,-13,5,-23,27,-1,5,9,19,16,-10,3,11,31,5,-16,19,-26,5,-7,28,35,-28,7,-17,9,-5,3,-1,45,26,24,31,-8,26,-4,32,5,-23,-14,-31,36,-1,-19,7,-4),
	(-1,41,-15,-5,-10,26,-9,-10,-20,-21,1,32,0,-36,-7,-8,-14,14,-4,8,6,17,20,-14,-17,31,20,5,-25,40,0,-4,21,12,5,7,-24,12,24,-5,-12,-38,19,22,35,3,23,18,-4,-4,-15,0,-15,3,4,-8,32,16,7,-19,32,-3,34,-25,-52,-23,-21,5,8,-4,-1,17,3,7,15,27,-11,-16,-20,-39,10,38,10,-27,32,-17,-6,5,0,32,14,25,-21,12,-17,-12,-9,13,8,-18,20,-15,31,25,-16,-14,-20,4,-23,-30,-2,29,-2,10,4,-20,19,-20,0,3,-7,-4,-10,18,19,9,10,28),
	(0,37,-28,-1,7,14,-30,31,-17,2,-5,22,-6,-13,-19,7,-17,24,25,-3,6,12,21,2,8,0,-23,-4,25,-16,17,5,-1,4,14,2,-9,7,-19,6,15,-12,-7,23,5,-9,7,34,17,14,-15,11,-21,35,5,0,14,4,10,-20,14,-8,25,-23,-42,9,-66,20,26,6,0,31,-10,-1,36,21,4,-4,-11,-27,-31,16,34,-26,19,-28,-30,5,-6,-7,-20,4,-31,10,20,-37,-21,-7,-17,20,14,-3,12,30,-21,-25,-18,-26,-18,0,-2,-2,-3,-14,-9,-12,8,-1,-14,11,9,4,-18,8,-13,24,0,13),
	(13,62,4,-1,-10,18,-6,42,-22,0,5,58,-22,-19,-42,14,0,17,-4,13,-2,-27,14,-6,12,0,-11,-21,18,-16,4,-11,-27,-3,0,24,13,-10,-1,10,0,4,-14,-3,19,-6,-1,36,27,-26,-18,-17,6,34,15,-22,-36,-9,10,17,4,-14,-2,-35,-26,-2,-78,16,26,2,-17,-6,-42,23,1,12,3,-5,-22,0,-39,4,16,-20,16,-42,1,6,1,18,-2,10,-14,13,22,-59,-20,-15,-27,15,6,-22,-36,-4,-30,-14,-15,-52,-18,-20,-5,-7,8,-12,-32,-29,-24,-19,-56,10,16,-14,1,-14,-25,-9,15,-10),
	(26,31,-1,-17,-2,7,-16,3,-6,8,-21,27,-28,-6,-51,0,21,7,-29,7,3,-33,14,-24,-40,15,8,-38,2,-57,5,-15,-3,6,-3,8,-19,2,-16,16,38,0,9,-21,3,-14,-29,-5,15,-4,11,-13,-3,15,15,-16,-26,-31,-15,-4,-48,3,26,-19,-7,-15,-98,-13,40,-26,10,-16,-89,2,-2,1,19,-42,-2,6,-38,-4,0,-45,23,-32,-13,2,-10,29,9,7,2,11,-9,-64,-10,-14,-39,-10,12,-20,-44,28,-38,13,-10,-31,-3,-4,3,10,26,9,-26,-31,-8,-11,-25,20,13,-6,-7,-37,9,-7,11,7),
	(37,15,-36,19,-40,25,24,9,19,-12,-27,35,0,-13,-27,6,-1,5,-39,-9,14,-36,33,-17,-5,0,-12,-24,6,-35,11,-12,-19,16,1,-12,10,23,-16,-12,20,-22,23,5,-22,-17,-4,28,-31,-13,41,16,17,-1,26,-26,-33,-10,-3,10,-46,-6,3,4,12,-36,-70,-5,14,-7,43,-6,-36,6,0,-3,0,-42,-41,-4,-14,9,19,-73,44,-41,-5,20,-2,-7,-1,1,-18,24,-6,-29,-10,-18,-32,-12,30,7,-41,22,-17,36,-40,-12,-5,-18,-4,-6,25,13,-9,27,4,30,-30,14,-16,18,-3,-43,-7,16,-9,-8),
	(36,12,-27,1,-26,13,5,8,30,2,-21,7,20,13,-28,-6,9,15,-37,-2,18,-46,-23,-31,-15,48,10,-10,-17,-15,20,-31,-7,-1,-9,2,-16,32,-35,-16,21,-29,10,21,-1,-34,5,44,-38,-12,44,-2,-4,12,29,14,-42,-9,-42,-12,-54,-13,35,-23,-1,-32,-31,-7,0,-6,33,-9,-28,-18,10,30,3,-32,-27,8,-17,-11,39,-84,34,-67,-21,19,15,-35,3,-12,0,-1,-18,2,9,-12,-33,-39,28,9,-32,25,-11,36,-40,-11,-38,-24,0,-23,20,-11,-20,0,0,0,-31,-3,-19,25,20,-33,13,5,-9,-60),
	(47,23,-1,15,-26,13,-8,-6,-4,-13,-23,16,16,19,-25,-11,-11,35,-27,-8,59,-13,-6,-13,7,10,42,-19,10,-40,3,-12,-32,-2,21,-4,0,5,-51,-19,0,-16,-16,7,-22,-40,-33,60,4,-34,-5,2,-3,33,24,7,-7,15,-36,12,-6,16,23,8,30,-31,-2,-36,-20,-23,-10,30,-2,0,5,-12,-13,-29,-20,-29,1,-5,10,-53,27,-59,12,9,-6,-32,37,2,6,-3,-4,-21,-6,-30,-3,-12,-4,22,-49,24,-6,16,-15,-12,-50,-32,5,-19,-35,-17,-21,-16,-62,14,-17,5,0,43,26,-24,2,5,-15,-37),
	(30,-24,9,34,19,34,4,11,32,-26,41,-25,34,37,-31,14,1,10,-57,-6,24,-31,-32,28,-4,21,4,11,29,-4,44,-10,-17,-16,35,3,5,30,-7,-41,-26,0,36,33,-61,-18,-23,40,-58,-37,-20,-12,-12,58,26,-14,0,-23,-61,0,7,21,27,-21,4,-56,27,-25,-7,-31,28,11,35,-32,13,10,2,-6,-44,-14,4,-25,13,-34,32,-5,32,41,-32,-18,0,-22,-5,71,-50,-19,-16,-15,11,-13,5,-16,-34,-7,7,0,-32,-14,-34,-12,-4,9,-24,-42,-56,-3,-33,39,10,-20,32,65,3,-27,33,-14,-7,2),
	(0,-55,2,1,-1,51,-9,9,45,-60,34,-36,34,4,-23,33,56,40,-38,15,0,-18,-15,-1,-7,42,-27,13,14,-17,35,-29,0,-30,21,-3,29,39,-4,-40,-47,-17,39,52,-15,11,5,-17,-41,-2,-30,3,-5,7,37,25,-10,-4,-23,-20,-6,40,37,32,31,-40,2,-25,28,-33,23,2,-1,22,-8,31,22,-3,12,-1,-20,14,31,17,22,-20,14,10,-9,4,-49,-14,7,11,2,6,-47,-2,-5,-29,27,-6,-41,0,-11,4,-16,-4,-3,-27,-9,28,-11,-7,11,2,-5,14,0,15,39,55,23,32,33,-18,25,1),
	(5,-9,-10,25,29,14,10,42,-4,-23,22,-31,25,12,-25,30,12,16,2,34,24,-11,19,6,-14,10,-10,33,27,-4,3,19,3,-14,31,-10,9,-8,-7,-22,-42,6,24,2,-6,-29,4,-5,-21,0,-4,28,-17,-23,21,5,-19,-5,4,-16,2,42,11,4,20,-11,-24,0,-16,-5,-22,-19,37,29,-31,6,2,-13,2,9,-19,0,-19,30,5,11,-16,-6,4,-23,-22,9,3,12,-16,-27,-28,-10,-36,12,43,0,-17,-30,2,6,-31,-27,19,-7,-35,9,-13,3,-20,7,1,44,10,17,6,3,24,-17,17,-4,27,25),
	(-18,-12,-19,9,15,6,-3,-3,-2,-13,2,8,3,-1,4,-14,-8,5,13,16,3,14,-12,-4,12,-1,-16,-4,-5,-14,7,18,13,-11,-1,4,-5,-1,11,10,-3,0,15,-8,-17,-16,19,-19,-14,-3,-14,-8,8,3,2,2,11,-10,14,10,19,6,7,7,8,11,12,9,12,-10,-7,-8,-8,-5,-15,4,-6,-6,-18,7,13,-1,-12,-6,-15,-3,-20,-11,17,18,13,-19,-1,11,-12,17,12,15,-11,16,3,-5,2,-19,0,-7,8,-10,7,20,-18,18,17,-15,1,-19,-8,13,-6,11,16,-10,-1,-15,-5,9,-3,11),
	(0,-20,2,-5,0,-5,-1,14,-13,-12,4,4,14,-1,3,4,-7,20,-4,21,-8,9,-7,27,4,-24,9,29,-7,26,-14,-8,29,-20,7,-17,-13,-11,-16,13,-10,-22,22,6,0,-15,-5,-20,25,-16,30,16,-2,8,13,4,2,0,17,-8,-5,10,-3,21,1,15,27,18,17,-18,-8,-3,1,27,12,-2,-16,14,-24,21,-9,15,-19,25,21,16,-26,-4,8,-6,14,27,-12,24,23,-2,25,-7,-9,21,-6,0,8,20,-11,18,-17,13,7,-11,9,-3,-9,3,11,27,1,-3,13,21,-29,-12,15,-2,7,1,13,-9),
	(-8,-3,-3,-10,6,5,10,9,5,-14,22,26,17,-29,-26,24,9,7,27,19,-17,-4,-8,-44,-2,31,-26,-10,6,-10,45,-11,0,4,3,-11,5,35,-9,-5,-12,24,-13,-20,18,-6,16,15,-5,-19,-21,31,22,3,-7,17,0,-32,-39,-12,-10,16,0,13,-44,-13,-37,3,-12,-4,7,-28,-22,-34,-34,9,25,-4,22,18,-15,12,35,-4,-25,2,15,-20,2,-28,5,-30,-25,-18,-19,3,0,25,4,-20,14,-2,-36,8,26,12,-28,-21,0,-8,5,44,-20,-5,8,-14,-14,30,3,-27,28,18,-26,-6,15,20,21,-7),
	(0,-21,-11,11,8,5,-22,13,23,-20,25,8,38,-65,-30,14,44,-24,34,33,-40,-29,0,-45,-48,39,-15,16,51,-17,0,-7,22,-5,0,17,-17,9,-4,21,5,-8,-19,-41,37,-1,9,-17,-17,-5,17,71,-34,26,27,0,-39,9,-38,0,-15,26,31,-24,-5,-43,-70,-12,-10,-1,-1,4,-57,-28,33,46,7,50,1,38,-25,42,42,17,-2,-12,7,38,-11,-25,-28,-6,-16,-15,-45,33,-24,15,17,-14,0,-14,-5,5,-13,5,-40,-26,41,0,-29,36,20,-9,-1,0,-10,35,-22,25,36,-22,-2,-64,54,14,29,-13),
	(-12,-21,-39,9,5,-4,-15,19,7,-33,17,-16,9,-48,-16,16,15,-10,-19,-1,-17,26,9,-48,0,16,-45,10,10,2,7,25,14,25,-13,36,-17,23,-1,6,8,-7,-15,-18,29,-18,-2,9,13,-12,14,36,-8,21,34,-26,-16,3,9,-5,3,10,12,3,-17,-14,-48,4,-2,8,18,26,-30,-19,-1,-5,-8,25,-11,18,-41,56,19,27,14,1,-8,-15,-39,-48,4,27,-27,-9,-56,48,-28,-1,23,-33,20,-36,-7,17,-33,0,-17,-24,28,20,-23,36,-10,13,2,5,-6,12,11,25,19,-2,10,-60,26,13,-17,6),
	(-23,-24,-38,22,-22,-7,17,-22,22,-25,-16,-5,2,-31,-6,1,0,13,-25,13,-11,34,-4,-26,32,22,-59,28,-45,-1,31,6,50,0,-11,-7,7,13,-6,-3,2,-10,-12,-65,19,-41,-21,7,-9,12,-2,16,14,35,28,8,19,9,9,3,10,-16,-21,5,-19,3,1,-19,-41,2,-11,-10,6,-16,23,-12,8,33,-33,10,0,57,10,-1,-4,-25,-1,0,-25,-16,-6,28,-24,-9,-28,44,-3,22,14,-7,-7,-34,0,11,-3,5,-12,-16,20,17,5,37,1,-10,-5,2,5,27,23,27,4,5,-36,-78,-26,4,23,16),
	(-22,-4,-66,19,6,14,-28,-29,14,-18,6,-20,19,-33,2,-6,-19,42,-2,15,-1,11,-3,3,3,0,-41,-6,-11,-5,36,36,-5,2,8,3,-23,4,-31,24,11,-18,-12,-48,-1,20,-11,-10,-7,21,31,32,10,7,23,10,13,-16,-14,-19,25,5,-6,-21,-70,4,42,-26,-48,-21,18,39,31,-20,31,0,17,19,-12,-19,-19,23,0,-5,30,-27,-10,30,-17,-4,1,-5,-14,-28,-54,17,-15,-19,44,14,-23,-27,29,15,0,19,-32,-22,-6,-21,-26,7,-14,20,-12,2,5,5,0,13,-4,11,-37,-64,-25,-4,4,-8),
	(-21,-13,-67,19,6,1,6,-38,32,-10,41,-15,27,-55,-16,12,14,13,15,14,-7,45,13,-13,-23,30,10,24,26,-7,9,19,-17,-2,5,8,-4,-10,0,8,6,14,-54,-49,15,5,4,-13,-3,11,36,22,-9,-4,1,-1,-26,15,-23,-14,19,15,29,18,-34,-4,-4,29,-75,10,24,12,10,-25,42,1,8,21,-5,20,-23,-11,33,10,-1,-28,-8,0,2,-8,1,0,-21,-1,-35,-1,27,-17,15,-6,14,-19,25,34,6,45,-45,-10,-19,-28,0,17,28,-12,-25,21,5,-1,8,-6,12,-2,-38,-71,-33,-27,4,-8),
	(-7,27,-82,17,2,20,18,-15,1,-14,46,-20,46,-42,-20,6,4,38,3,24,9,11,30,0,6,24,6,-2,-13,26,29,0,9,-14,2,-6,22,-8,-39,21,23,-3,-72,-40,-10,-17,2,-26,-7,-23,17,28,36,-2,14,-32,0,8,-7,-5,5,-2,11,-3,-58,-14,37,-2,-76,4,3,16,20,0,19,-8,3,-4,4,12,-20,8,11,-6,6,-44,-8,21,-16,11,0,-5,3,3,-27,-39,22,2,16,16,25,-8,0,25,4,23,-16,-20,-16,-12,0,12,18,1,9,6,-7,26,-7,12,-2,12,-43,-73,-11,-12,24,1),
	(-20,20,-81,6,-25,19,35,-15,3,-2,28,-17,48,-29,-65,3,-9,16,2,17,-15,-28,8,-12,0,-4,36,2,-12,-2,-9,13,2,20,30,-29,-8,20,-17,22,23,4,-51,12,0,-34,-6,-28,3,2,0,15,23,-22,15,-23,3,-3,-8,15,11,36,14,-3,-41,-1,24,31,-67,-4,-2,20,17,-20,31,19,0,6,0,18,15,-15,-1,-19,-7,-8,-34,0,-20,5,-17,3,-21,20,-11,-24,20,-2,36,-15,26,3,6,15,18,13,-50,-20,-36,-31,-9,4,0,0,-27,21,26,-5,-32,0,12,25,-22,-61,-14,-9,12,-18),
	(-4,12,-87,-14,-17,13,21,10,3,17,28,13,43,-4,-83,-5,6,18,30,-6,-22,-17,44,5,-6,20,37,0,-16,-18,-6,-28,-6,28,39,-10,22,14,-40,-24,11,35,-15,42,17,-42,41,6,-18,4,-6,0,6,-30,12,-43,-17,11,23,7,12,35,22,-20,-43,21,32,31,-84,1,13,-18,22,-11,19,11,2,4,-31,5,-5,3,-18,-8,5,-40,-27,34,-11,-1,-41,-16,-11,27,12,-11,-1,-6,2,4,21,33,29,-19,9,31,-18,9,-24,-28,-9,21,33,0,-8,21,20,0,-36,7,-6,42,-7,-16,8,18,-3,-22),
	(0,10,-43,8,-3,12,-22,22,-29,27,36,-4,2,30,-30,30,2,10,19,24,-13,-32,57,17,-11,-3,22,-18,-43,15,14,-18,18,16,23,-12,26,23,-35,-12,14,-8,23,23,-9,-16,28,-6,-10,-18,-21,7,8,-52,45,-44,-23,-13,-8,-3,-9,40,12,-10,-30,-1,15,33,-89,11,-6,5,37,-22,1,7,14,-10,-14,22,-2,0,-29,-22,16,-13,-22,10,10,-1,-8,-2,8,28,13,-26,14,-28,9,18,22,24,-18,10,9,22,-45,4,-25,8,-28,35,31,6,-50,26,4,40,-29,19,2,23,21,40,0,5,26,-12),
	(-4,1,-37,-1,1,24,1,26,-22,42,28,-4,3,28,13,17,-7,12,8,4,-24,-69,30,10,19,0,-13,-7,-15,19,-25,-13,-4,19,33,-36,6,6,-47,-17,25,-4,32,11,4,13,22,-6,1,-20,14,14,15,-51,9,-15,-26,-11,13,-12,-2,25,12,-20,-17,11,21,1,-74,14,-24,-1,16,-25,-23,15,12,11,8,0,21,-5,-35,9,19,9,-39,40,-17,-12,-7,-6,31,25,-22,-22,-17,-12,8,28,-8,40,-4,10,7,8,-16,-3,-31,-24,-15,22,18,-32,-25,7,7,19,-15,26,20,3,56,38,-15,24,32,-1),
	(-11,-14,18,-18,-24,-14,0,18,-5,39,21,-7,-2,-8,0,5,11,16,15,24,7,-51,4,-24,21,-20,-13,12,6,9,7,24,27,-11,4,-8,-7,14,-42,9,-4,-9,17,-1,-15,27,-6,30,7,3,13,1,-20,-14,5,-12,-7,-3,-7,3,10,26,11,-24,-5,13,39,22,-44,-14,14,16,35,-10,-1,10,-6,-9,-12,7,-2,-16,-22,2,6,5,-34,28,-6,15,9,-7,29,9,-14,8,18,-9,4,25,-14,36,20,18,-5,-4,-35,-13,-39,-10,5,4,7,-9,6,16,25,20,4,6,29,-38,21,24,-17,14,-2,7),
	(-26,1,5,18,5,10,3,9,-39,7,27,-39,-9,-57,18,22,12,-9,7,-2,-15,-79,-12,-29,-26,-10,-20,-8,33,30,-24,14,13,3,-14,-32,-1,10,0,10,51,5,49,2,-12,17,-7,7,-16,11,9,0,-36,-6,4,-27,0,3,-7,15,-12,11,-6,-28,1,8,38,15,-49,-18,11,5,15,23,10,28,-14,-3,-10,8,20,-16,-27,9,14,30,-13,19,2,4,40,-1,-7,14,-21,3,-11,-18,21,5,7,-3,-13,6,-19,-2,7,-3,-36,-17,0,18,9,0,-5,27,21,31,-7,24,0,-16,-4,32,1,7,25,17),
	(-22,0,-11,-4,12,-1,-30,-14,-28,-15,9,-24,27,-66,16,2,2,2,3,6,0,-58,4,-7,-20,28,-22,10,5,26,7,24,0,21,15,4,0,7,10,-1,22,10,26,-3,-8,18,19,16,12,-5,-10,2,-38,-8,-12,-15,17,0,-4,2,4,1,7,9,-32,-9,18,39,15,17,30,24,-15,-19,20,-3,3,5,-15,-9,19,9,-12,-15,-3,-12,34,21,-15,0,37,6,26,-3,-23,25,2,-20,29,-6,-5,9,21,32,-42,22,-22,19,-6,9,-4,37,8,1,19,-13,18,29,-7,3,21,-9,2,38,-22,-10,-2,-7),
	(-9,10,2,8,16,1,-31,-31,-21,15,22,-24,23,-48,34,26,13,-1,-7,15,-25,19,0,-23,-20,1,-13,-4,6,28,20,15,10,23,13,0,4,41,-1,-6,21,-19,18,-3,0,-9,10,16,3,9,-24,9,-32,-6,0,13,0,6,-28,14,-13,20,-22,-26,-35,-10,-6,-2,5,-10,-6,14,-15,11,1,-9,-6,11,-6,1,22,-2,4,-22,30,8,18,7,-3,0,32,2,3,-6,8,-4,23,-18,14,-10,19,-7,28,24,-7,-23,19,10,21,-18,8,44,-14,14,1,-14,2,14,29,20,-16,8,0,26,5,5,9,3),
	(29,51,34,-1,-5,0,-16,-38,-2,0,34,16,20,-48,7,-2,1,18,6,9,-11,44,39,-30,2,10,-16,-6,-8,17,34,18,-14,22,9,29,-21,30,4,20,17,-36,21,-19,7,0,-9,35,-15,-24,-24,7,-19,3,10,6,17,9,-20,6,29,11,1,-3,-38,-7,-1,11,-21,2,26,18,-26,-17,16,7,6,-15,-23,-17,29,5,-3,-8,46,-15,-6,8,-1,-21,29,19,17,-17,-14,-9,-12,-26,0,-1,-10,-5,40,44,-28,3,2,5,7,-23,11,41,11,-3,31,3,-3,-4,8,-3,13,4,-20,42,2,-16,-5,7),
	(24,45,-22,12,30,27,-30,0,-30,0,41,1,4,-34,-38,-2,29,33,-9,11,-14,9,25,-11,-6,5,18,-4,5,22,1,-2,-20,41,25,28,-20,11,-2,22,20,-24,-5,17,26,13,6,19,-4,1,-37,-1,-15,33,-9,-10,12,-32,-32,17,16,-10,-4,1,-54,-11,-53,27,19,1,25,0,-19,8,31,7,-13,-11,-22,-34,0,25,23,-37,37,-12,0,-1,17,25,0,-5,4,-9,-20,-30,16,-7,24,-6,1,0,27,31,-19,0,-2,-2,-6,-14,-11,32,3,-7,-8,-14,21,6,-4,4,-6,4,-12,22,3,-3,-22,18),
	(47,50,6,11,-26,6,-10,11,14,-2,9,22,7,-38,-9,-5,-3,16,20,-13,2,-10,28,-15,0,15,-14,-5,-15,15,23,-20,-23,36,17,22,-19,-23,10,22,3,3,17,17,-6,-7,-8,18,-8,-14,-19,-20,-14,35,5,-3,1,-15,-17,-18,3,27,14,4,-36,0,-119,-3,22,16,38,33,-35,5,35,-6,4,-8,-13,-28,-16,-15,11,-41,34,-23,5,10,-9,-4,17,24,-29,3,-14,-44,5,-6,-19,-2,16,5,-17,20,-13,-1,3,-36,-6,-1,-15,26,23,-7,-12,4,-21,-6,-12,16,20,-5,-21,31,-34,1,-20,6),
	(23,19,3,-3,12,17,-26,10,15,-5,-1,42,3,-15,-53,-15,3,15,-1,23,5,-32,24,-10,-10,6,-14,4,18,-5,15,-5,0,-9,-17,30,-24,21,3,5,4,-17,-11,16,21,-28,0,42,10,-2,-14,9,-10,22,26,-27,-42,-33,-18,-9,-38,7,12,-12,-24,-16,-107,-9,20,-8,28,12,-57,7,37,4,-3,-16,-32,-1,-11,0,6,-58,34,-42,-18,-10,12,4,-5,9,-29,27,14,-37,9,-19,1,-6,4,-10,-11,25,-18,-5,-23,-52,-22,-26,-3,4,19,6,-28,-12,1,-20,-55,5,-3,0,-22,12,-22,0,-9,-5),
	(28,4,-7,5,20,39,-10,35,20,-14,-1,39,0,-7,-42,-5,12,22,-12,4,-30,-27,26,-39,-25,34,-4,-1,16,-22,5,-18,8,16,6,11,-5,-7,-8,-1,-8,-19,0,-7,11,-8,-48,22,0,-35,2,7,2,14,-4,-18,-41,-17,6,-9,-57,8,-11,9,16,-6,-69,1,18,-18,17,25,-67,-2,30,5,-1,-17,-38,22,-28,11,-8,-17,22,-42,-19,12,15,16,15,-12,6,12,-2,-64,-39,-15,-52,8,19,-3,-33,9,-9,19,-7,-40,-25,-36,-12,14,7,8,22,-14,-28,8,-60,26,22,-4,-9,17,-25,12,-6,5),
	(43,31,-29,24,-4,26,0,26,-1,13,-16,13,32,5,-71,11,-5,30,-42,21,8,-17,4,-37,-5,29,27,14,-15,-27,-3,-43,-23,23,0,-15,-9,12,3,-24,36,1,-14,11,2,-33,-25,33,0,-10,21,14,-26,25,18,-7,-36,-46,-10,-9,-69,-18,17,3,6,-11,-35,-9,-13,-26,35,-13,-56,10,26,-4,18,-25,-51,-29,-4,10,-7,-19,27,-50,10,15,18,-28,-25,-13,-19,11,-15,-12,-1,11,-44,-8,27,0,-45,28,-25,4,-8,-24,-19,-42,2,12,15,-3,-3,3,-38,0,-18,15,25,19,-36,-23,-29,21,-6,-21),
	(38,16,21,33,-17,15,5,22,36,-1,17,5,27,17,-26,-3,-38,5,-2,-2,6,-57,-6,-14,0,52,29,16,6,-45,29,-14,6,-5,13,8,0,5,-18,-6,9,-26,-3,-7,0,-17,-28,-2,-38,-28,-15,-20,-27,42,10,9,-42,-3,-41,-1,-35,3,16,-2,27,-36,-39,-30,-8,-19,19,10,-37,-8,15,3,5,-20,-35,-5,-26,-2,-6,-34,32,-14,4,34,22,-17,13,-21,-16,-21,-6,-24,22,9,-42,-6,20,0,-57,5,-26,16,-4,-13,-26,-40,-2,-13,3,-22,25,-3,-38,-8,-17,-4,1,3,-25,7,-14,-8,-20,-19),
	(79,21,15,-7,-7,-1,11,-37,-9,-16,-7,-19,34,40,12,-11,-4,6,-23,-19,55,-47,-24,18,6,5,-21,-1,8,-33,12,-12,-4,19,-7,-1,12,-2,-40,-21,29,-35,-4,19,-15,-3,-46,34,-47,-13,-3,-3,-3,67,12,14,-34,-4,-27,-7,-29,4,16,-2,42,-29,0,-24,-12,-39,21,8,19,10,0,3,-2,-8,-10,-9,-15,2,22,-65,28,-25,-3,24,-16,-27,23,-15,-29,5,36,16,26,11,9,-9,-13,-23,-20,-1,1,-1,3,0,-50,-13,5,7,-34,-15,-22,-7,-25,-27,-44,-30,-1,3,29,40,22,38,-27,-29),
	(33,33,35,-8,2,-3,-3,-26,-9,-28,22,3,25,56,-29,1,3,40,5,-9,53,-37,-25,4,17,32,-27,-18,12,-22,59,12,-30,-11,17,-8,19,31,-29,-28,-33,-14,-8,11,-41,11,-34,13,-51,-36,-52,-35,-11,44,-5,-26,-7,-12,-64,10,-2,8,2,-2,16,-9,12,-2,3,-29,10,7,14,-4,22,-28,-4,-14,-42,-31,28,1,7,-66,25,-30,12,19,-2,-12,-19,-29,29,12,-39,18,-2,30,3,-25,8,14,5,6,7,-12,5,-10,-11,-41,2,48,-4,-28,-38,-3,-16,12,0,-22,16,30,4,5,0,44,8,-2),
	(-14,-47,-24,9,16,46,-3,3,20,-7,26,-29,25,-1,-23,-9,36,10,-39,0,-8,-20,22,0,-15,13,4,1,21,19,7,9,-19,-7,5,25,2,21,-29,-9,-23,5,15,35,-2,30,-31,19,-19,-27,-8,0,-16,7,27,1,9,-15,-13,0,-11,7,27,17,34,-36,37,-12,9,-21,35,32,5,9,-4,13,-3,-2,0,-14,-5,-16,15,0,28,-10,-4,13,-35,4,0,-30,-23,29,-42,-23,-23,-17,31,12,-15,0,-31,-21,-8,0,8,4,0,-2,-23,22,-1,-12,8,-14,-1,5,11,-8,-10,15,-10,33,19,-8,3,24),
	(2,18,8,17,15,-5,-15,16,-10,-2,6,7,4,-4,9,-11,-3,10,-15,-13,0,9,0,-16,-13,0,5,7,-8,3,-6,-7,-3,7,3,21,12,14,16,18,15,15,17,24,-17,-12,16,11,7,-12,11,-24,-21,-11,7,-11,20,-9,9,-9,11,14,-21,-17,24,6,9,0,16,11,-8,18,-6,-17,5,-17,-18,-2,-8,-23,-6,-19,16,-2,18,20,12,-12,1,12,16,-19,-21,-2,-2,7,5,14,1,3,3,-4,4,-11,0,-19,2,-7,-12,7,-12,-2,-7,-21,6,-21,6,13,6,-4,-15,22,9,-5,-13,-8,3,2),
	(-5,14,13,-12,-10,-2,-3,15,16,2,1,-19,-12,7,-21,-6,-11,21,-20,-4,-2,10,19,-10,1,13,-13,-12,17,22,12,20,-20,13,20,-12,-7,11,-10,2,-9,-7,19,8,-24,-5,20,-14,-25,12,13,0,-10,0,-10,9,-9,-25,11,15,11,19,17,19,-7,5,-16,-17,-5,-10,0,18,0,-15,23,11,11,1,8,-13,5,6,-16,15,-11,-13,-3,14,-6,24,0,9,-19,26,-26,-13,18,2,-12,14,-21,-3,11,-11,21,4,17,-2,23,0,4,-10,-22,-14,4,4,-4,-4,-1,-7,-21,21,-10,-15,-11,-11,-7,-13),
	(15,-18,13,16,-5,-9,-9,19,27,20,9,-10,0,17,11,10,-7,-8,2,-3,-4,0,29,-39,-7,25,3,9,21,-20,10,21,-15,-37,13,-7,12,-15,7,10,0,12,-10,-8,3,14,19,-12,-19,4,6,-18,-4,-6,0,6,-35,8,15,-17,17,31,19,-4,-12,-15,-9,12,21,10,18,15,-34,18,-17,11,-7,19,-9,23,-24,1,20,10,3,-21,-28,15,-8,-6,12,17,0,5,-18,10,28,30,-11,13,-14,6,13,16,-24,19,12,-17,2,-1,0,0,-10,19,5,3,16,-1,13,5,-25,-9,-14,-10,23,-19,1,-13),
	(-9,-9,-14,32,-23,5,13,38,40,-28,39,-1,15,-39,1,14,52,0,30,52,-19,-8,14,-5,-46,16,-9,53,11,-21,10,-21,9,-21,8,-1,-15,20,17,-32,-23,-46,0,-5,9,6,18,-6,-20,-25,6,33,-27,3,18,7,-16,5,-33,10,-35,31,21,1,9,-12,-15,0,3,-3,11,1,-8,0,-24,12,-4,34,17,47,6,16,36,-18,20,-40,-9,-11,22,-9,14,-13,-23,10,-53,15,46,1,-44,-39,8,12,10,1,0,13,-21,-46,17,12,-25,29,12,-8,32,36,1,6,20,-10,44,15,-14,-7,25,-3,23,-36),
	(-30,-42,-34,43,18,29,-1,25,40,-36,40,-16,14,-27,-23,21,67,27,30,35,-38,-6,20,-38,-25,23,-35,36,22,4,0,-10,12,2,-25,-2,-42,31,0,-15,5,0,-21,-29,20,-7,43,-8,-11,-15,20,27,-25,1,26,-12,-14,11,-26,-3,-4,39,55,15,-1,-20,-34,10,5,-21,33,15,-39,1,4,1,3,46,-38,27,8,22,50,3,48,-11,-6,-2,-24,-9,-33,-8,-17,2,-23,8,4,13,-12,-44,16,4,22,46,-37,24,-36,-12,41,-7,-38,9,-13,-15,-4,40,3,-3,-4,10,15,16,1,-52,7,-5,8,0),
	(15,-34,-40,11,33,-1,-33,12,16,-7,31,6,23,-21,-30,2,-6,15,-1,2,7,0,17,-49,-13,-5,-38,-3,2,19,29,-5,6,25,-24,8,3,10,19,4,27,23,-5,-27,8,-27,-14,0,3,-6,-17,31,0,6,5,-1,1,13,-10,-1,-14,-6,-11,-25,18,-15,-6,19,-10,-11,27,-1,-26,-18,19,-6,9,21,-8,-10,-16,3,8,17,19,-12,-13,3,-12,-21,16,-8,-63,18,-26,27,-11,23,-24,-29,24,-18,0,5,-29,-3,0,-12,31,15,-11,19,-20,4,12,1,-26,2,-5,24,0,27,-1,-72,7,-4,-19,17),
	(8,-25,-57,13,18,7,7,-9,20,-8,26,-22,19,-12,-8,-14,-13,16,-20,8,12,31,14,-19,19,-6,-9,7,-11,4,40,1,0,-8,1,31,2,-7,28,-6,24,7,-35,-73,7,7,-27,-17,-26,4,14,5,-4,12,-16,15,20,9,-4,-18,-18,4,6,2,-46,3,6,-35,11,-27,-13,0,-27,-34,27,-4,-6,-17,-7,3,0,-1,-2,24,15,-32,-1,-7,0,-7,-17,-16,-13,-10,-20,20,-11,-13,-3,-37,-9,-6,-28,19,-25,7,16,-5,45,25,5,13,-36,-29,-14,-14,-34,16,16,1,-13,9,-43,-78,-18,-6,17,21),
	(-11,-11,-47,3,26,-19,15,1,11,-4,6,-15,-9,-52,-13,-11,-35,9,3,6,19,60,18,-11,-8,19,-14,16,-16,-12,27,26,7,5,14,7,-4,20,7,7,29,-12,-62,-47,5,-19,-14,-13,8,7,27,14,-2,17,18,-24,28,-17,8,-14,22,-11,-11,22,-69,-22,24,-25,-3,-1,14,12,-23,-41,27,3,16,-11,-31,-18,-26,7,-19,30,50,-57,-10,-17,-18,-29,4,27,8,-6,-54,23,-15,0,-23,-12,-4,-6,-9,39,7,36,18,-8,40,-33,3,40,-10,26,-6,24,-11,20,27,-1,-3,7,-44,-59,-30,2,5,12),
	(-24,-19,-42,12,-5,0,0,-12,31,-32,21,-7,20,-37,-35,8,-20,33,0,16,-21,46,6,-3,-2,26,-1,-14,10,2,2,28,15,-14,-4,13,-21,-3,11,-20,39,0,-36,-37,24,3,-12,7,-7,-3,13,0,31,-7,13,-21,-11,-9,5,-17,30,-11,-3,-7,-66,-24,19,10,-13,-2,37,3,4,-3,9,23,-8,0,-33,-12,0,-23,-12,6,34,-38,14,-7,-23,-6,-19,9,-13,-12,-37,32,35,7,-12,-8,5,11,13,51,-15,19,-7,-3,37,-22,-2,2,1,6,11,5,-13,28,41,37,-22,0,-59,-53,-18,-21,-2,9),
	(-13,-29,-61,8,23,25,24,-10,36,-14,17,0,12,-33,-21,14,-4,7,-7,13,-9,21,34,-9,0,8,19,0,8,26,15,27,0,13,5,4,-24,-23,22,11,17,22,-56,-24,16,-1,-24,16,-12,18,18,7,7,-9,16,0,-3,5,-10,15,5,-24,-17,4,-49,14,-7,36,-47,4,6,18,10,-14,37,24,-10,-7,-13,-2,-2,-9,30,-16,5,-8,2,16,-9,-21,7,-12,-21,11,-25,12,2,-6,17,21,0,-4,28,13,-14,7,-27,7,21,15,-9,40,16,9,-8,34,5,25,18,30,-15,8,-20,-34,-14,9,0,-5),
	(-15,-34,-41,-3,18,3,30,11,25,3,38,7,14,-28,-53,14,-13,32,5,-1,-4,1,7,-3,16,-4,-9,-9,-5,-2,-8,-10,5,-3,20,-29,-12,-9,-6,-3,29,10,-36,-6,-5,-40,5,0,-4,8,9,-6,5,-6,2,-14,-16,-21,7,7,5,-14,3,-4,-20,-1,14,45,-68,-3,-6,-7,4,-31,32,1,5,-1,23,10,5,-6,-14,-15,7,-3,9,3,-17,13,7,4,-19,-4,14,-8,-12,-5,0,25,4,11,20,3,-6,6,-34,-25,30,14,-20,22,10,-23,-9,-6,17,7,2,2,-8,34,14,-10,-9,7,3,-27),
	(12,-1,-31,9,8,-2,20,-27,27,7,17,-15,10,8,-43,32,5,17,-12,0,-45,-22,33,19,-14,7,14,-3,-18,8,-4,-8,-14,15,0,-16,5,11,-18,7,25,11,-44,31,-18,-14,4,26,-10,6,16,-7,9,2,9,-24,-26,12,13,-8,10,-1,21,-8,15,27,20,30,-23,34,9,-15,10,-8,19,22,-6,-6,-6,4,10,-30,3,7,-13,-34,16,6,-4,-13,-30,0,-12,23,15,11,-1,-19,0,18,-6,-3,18,13,25,1,-8,-7,-6,5,-16,34,11,-23,-31,34,22,28,-18,-3,34,15,-5,26,-8,5,2,-14),
	(-4,23,-16,-28,22,7,15,22,-7,23,9,-25,-8,-19,-25,16,1,18,11,18,-31,-39,26,30,-6,2,-2,-24,-15,13,10,-19,-2,8,12,-20,17,11,-9,8,37,14,-16,24,24,-32,2,-16,13,9,1,-8,11,-9,30,0,-28,10,-6,-2,-1,10,11,-19,-5,13,37,27,-48,29,-5,18,11,-14,-9,31,19,8,14,-2,12,-14,-38,-3,17,-17,0,29,-3,0,-29,10,19,35,12,2,-11,-22,0,11,-1,37,10,-7,5,9,-33,7,8,-14,1,21,18,-7,15,-7,22,39,-18,32,18,29,18,32,-39,3,39,-26),
	(10,0,-27,0,-9,-6,2,-25,-26,0,31,-17,-20,-15,4,23,15,16,12,18,1,-73,15,-1,22,8,0,13,-11,12,-9,-12,11,18,28,0,20,2,-27,-9,19,19,11,21,12,6,-10,21,2,-5,0,-16,-7,6,27,-19,-29,-14,-9,-6,37,-5,-7,2,7,33,8,35,-27,11,-13,17,34,11,20,24,-1,17,4,23,-10,-1,-50,0,-6,12,6,7,9,-13,-5,10,-1,8,-33,-5,-7,-23,26,18,0,31,24,-21,-2,13,-25,13,-14,12,-23,38,28,-6,4,2,-6,32,-21,11,37,11,15,23,-14,13,33,-33),
	(-1,-5,-17,-15,10,-3,-5,-14,-5,11,17,4,-13,-45,18,49,-6,24,-11,16,-20,-84,-13,-15,0,4,-10,14,-1,2,-4,6,2,10,28,9,0,-4,-46,-3,37,-11,8,11,-7,-6,26,40,5,-9,2,9,-2,-9,0,-10,-26,0,3,4,21,-1,6,5,-3,-4,14,39,-23,-18,0,11,-1,13,-10,27,-16,0,0,-6,0,6,-36,-11,-3,0,29,13,16,-26,-6,1,9,5,-3,1,0,-11,14,5,-9,16,31,26,-16,-1,-19,6,-31,22,-32,26,28,-4,-1,17,8,48,-5,26,38,-4,23,22,-38,20,14,-3),
	(20,-16,10,-6,1,26,-31,-14,-5,3,29,-21,-17,-28,27,35,-2,0,16,3,-25,-60,17,-25,-14,25,-27,3,0,20,-29,9,3,18,16,-9,-20,8,-35,12,26,8,47,-3,10,17,-2,33,-6,-11,-21,-34,2,-6,2,2,-14,9,8,-19,13,8,-23,-19,-31,-24,36,42,-22,6,30,-7,-1,1,25,-12,7,-1,-10,-2,-2,5,-36,-3,45,-4,-7,4,-13,-19,23,5,36,13,-18,12,5,-12,47,-25,23,22,13,1,-30,13,8,34,-24,-19,-9,20,18,11,0,30,9,8,-23,19,35,-33,-8,51,-62,15,28,5),
	(-1,-1,8,-5,-5,17,-29,17,-15,3,29,21,-7,-39,21,25,0,25,-5,-3,-18,-30,6,-31,-9,-13,-21,-9,12,36,-22,42,-16,14,11,21,-16,14,-11,-13,43,-1,24,2,-6,26,-13,9,22,0,-23,14,-10,-13,8,-15,24,14,6,0,18,8,-18,-3,-8,9,2,50,-4,4,14,-7,-1,12,0,-32,-16,-4,0,1,-2,7,-20,-13,24,-28,36,21,-3,4,38,0,4,-8,0,13,10,9,13,-32,8,8,19,30,-2,-6,11,4,-15,-20,1,43,37,-2,-3,-9,5,10,-1,23,20,3,-3,31,-17,24,22,-9),
	(-4,6,7,19,10,0,-35,-15,-16,1,22,17,24,-41,22,34,-13,1,-27,5,0,18,7,-22,-20,15,-14,14,4,4,12,5,-13,20,0,29,14,16,1,0,25,-27,5,-12,3,0,-7,-14,-12,6,-22,1,-18,0,-20,-12,19,17,-6,-3,0,16,-2,-25,-13,-6,-33,17,1,0,21,16,-17,4,9,-39,-9,2,-15,-18,19,24,-32,-29,-4,6,26,14,24,18,29,10,1,-28,23,-18,20,-16,22,-42,0,13,32,-1,-23,-2,-15,5,17,-23,-2,53,22,12,8,4,-9,5,18,15,0,19,-4,20,-28,-3,-6,15),
	(37,15,-23,6,28,18,-10,-18,-9,-4,13,31,21,-32,13,6,19,-7,-12,-9,4,17,12,-11,-28,9,6,25,1,18,-4,-7,7,0,-7,30,-20,22,5,6,9,-20,-28,-1,30,-19,14,21,-2,8,-6,15,-24,-4,-1,0,27,6,0,-20,13,17,-21,-18,-48,-20,-23,25,-8,-4,4,20,-16,-20,29,-35,-3,13,6,-32,10,21,-15,-33,32,-47,8,5,31,-9,22,-8,23,-23,21,-18,12,10,3,-19,26,10,16,21,-7,-13,-13,-15,8,-29,-8,42,20,7,0,17,-9,3,7,7,11,-13,-14,42,-27,3,8,11),
	(22,38,-24,23,-3,25,-19,14,-9,15,40,9,19,-31,0,31,15,0,-4,15,-39,17,-2,-33,-13,7,4,0,2,-8,15,12,-1,32,-10,13,-16,25,2,10,21,-14,0,-1,0,-7,-14,31,-21,-23,-23,-23,-12,5,-12,-11,-4,-15,-8,-11,0,-1,11,-14,-22,-17,-71,38,-7,-10,39,2,3,-19,23,-15,21,16,-12,-23,-12,10,-12,-78,25,-20,-11,0,9,22,14,-9,-17,2,-25,-54,-22,11,-10,2,-4,19,-22,20,-31,-10,-21,-2,16,-16,-1,37,33,-27,-27,24,9,9,-5,37,32,-2,-3,54,-3,-4,2,23),
	(44,32,-19,30,9,42,-30,-6,-18,13,56,15,10,-22,0,1,31,37,2,26,-5,12,15,-16,-32,26,-6,-1,4,-15,10,6,-13,-6,4,27,-33,-3,-18,22,18,7,-9,4,28,-7,-16,1,11,-19,-31,-4,-26,25,1,-22,-26,-4,-32,-16,-23,18,-8,-8,-30,-38,-118,24,-7,14,21,5,-39,-12,44,-29,4,32,-28,5,-14,1,-3,-76,12,-45,-5,16,-19,20,8,-6,-28,0,7,-53,9,8,-34,-10,-4,7,-38,0,-24,4,-18,-16,0,-29,-11,39,30,-2,-2,0,-3,-15,-52,17,3,-8,16,25,-41,-10,7,-19),
	(43,43,-22,3,28,23,-47,4,12,-4,22,49,15,4,-25,3,22,9,-21,-7,12,-39,23,-8,-26,0,8,-8,-16,-8,13,-14,-8,0,-9,18,-31,-5,3,11,25,-6,3,10,20,-41,-33,11,-2,-28,9,7,4,36,10,9,-28,-41,-26,-13,-52,33,11,-26,-10,0,-86,15,7,-14,17,8,-84,-17,43,-27,-14,-7,-25,-15,-21,-9,-5,-33,15,-42,9,-4,-5,-10,-3,-17,4,5,-15,-65,-21,-15,-13,4,-4,20,-31,41,-14,-25,-16,-20,7,-28,4,17,10,1,0,-35,-32,-20,-45,3,8,-9,-18,7,-39,23,-5,9),
	(34,8,2,-1,29,10,5,35,-8,0,5,31,20,30,-27,28,20,6,-34,6,-2,-20,-4,-35,-43,13,-1,-4,13,-26,18,-26,-25,21,21,-15,2,24,-10,-21,33,0,-23,-9,21,-43,-64,16,10,-8,4,21,-37,32,11,0,-27,-50,-7,-8,-62,21,-4,-14,17,-30,-75,-37,-11,-20,2,-17,-84,-15,8,-2,11,-2,-13,-11,-30,-7,19,-30,13,-11,-3,15,-22,-23,-15,-47,-1,-2,-32,-42,-28,-10,-69,-3,6,-4,-41,0,-16,-2,-8,-59,-6,-34,-6,0,-10,6,2,-25,-40,19,-19,3,3,-14,-6,-5,-32,-7,10,10),
	(21,9,13,10,16,16,0,30,10,12,25,8,21,2,-35,9,-9,9,-6,36,-13,-39,-2,-13,-32,7,23,27,9,-6,31,-33,5,-9,4,2,8,34,-28,-27,0,-13,-13,-5,41,-28,-53,28,7,-16,-16,12,-14,-8,-25,3,-37,-35,-30,-6,-67,0,24,5,0,9,-20,11,-15,3,5,-2,-45,-9,14,-6,18,-27,-7,1,-28,20,26,-28,12,-25,7,13,27,-18,15,-6,16,-23,-26,-21,-16,10,-44,5,18,18,-81,7,-29,-4,9,-33,-32,-19,-14,12,36,4,32,2,-12,28,-32,9,20,-6,-25,0,-45,1,4,-24),
	(52,-26,-1,32,-6,16,16,52,14,-13,13,8,41,0,-8,36,8,25,-12,26,-4,-69,-13,-25,-9,20,31,2,9,-25,55,-36,-15,9,-16,-39,0,16,-9,-34,32,-21,1,15,19,-18,-67,22,-7,-37,-4,2,-35,18,-5,31,-37,-37,-37,-4,-37,3,-4,-14,24,2,-15,-21,-24,-30,0,-13,-18,-29,-27,12,39,13,-15,10,-3,2,7,-33,-5,-3,24,0,22,-58,-5,-18,-9,-28,-4,12,29,-5,-45,-14,36,-12,-32,27,0,-18,-20,-40,-15,-27,-7,26,-1,-44,-8,-28,-47,32,-24,-11,22,-3,-19,15,-13,6,-1,-24),
	(21,24,17,25,18,-2,13,-34,-33,-29,39,-23,70,38,8,15,-12,3,-51,-16,27,-7,10,-9,-6,13,4,19,3,-36,54,-18,-16,3,26,-10,-7,30,-16,1,1,-21,-11,9,-14,8,-47,-19,-19,-49,-34,-20,-21,65,39,12,-25,-18,-12,12,-48,52,7,-24,42,-16,-20,-38,12,-14,-9,16,-8,-11,3,-5,9,-7,20,-22,18,0,12,-10,26,-1,32,-5,-31,-30,-6,-23,-25,-9,26,-14,-4,15,24,-32,-9,-28,-27,-8,-4,-9,14,-13,-38,-11,2,55,-68,-27,11,-29,-61,6,0,-13,18,33,35,34,21,-3,15,-14),
	(35,-3,35,0,18,-8,-10,-14,15,-41,22,-4,21,32,-18,12,-15,15,-6,21,57,-3,-15,-2,5,9,-17,-7,19,-24,38,12,-7,17,24,0,13,40,-29,-20,-11,-41,-4,-14,-6,-22,-14,31,-11,-20,-10,15,-15,40,26,-5,-10,-18,-46,-1,-22,5,4,-38,4,11,11,0,46,2,-5,0,-1,-8,0,-9,-8,33,-15,-8,3,7,-17,-50,14,14,-9,13,-47,17,21,-18,24,-10,-35,19,-14,-34,-18,0,5,13,-14,7,-13,-35,5,-28,11,-36,0,20,-20,-57,-21,-21,-15,-2,-2,-2,27,35,-12,22,-13,30,32,-16),
	(-29,10,-36,12,44,-35,7,-19,-15,25,31,-4,-17,-25,-15,36,41,14,-42,20,-42,-19,31,6,29,-39,-10,-5,13,-11,-28,-39,33,12,9,7,31,35,-14,-5,-18,-18,9,44,-19,-11,13,26,10,-59,0,47,3,-9,-17,-20,-25,17,13,-19,-2,38,21,-23,36,1,37,29,16,5,-24,-5,-21,13,-34,30,-31,-13,-32,35,29,-23,15,0,3,51,19,33,-45,-19,25,-11,21,50,-57,1,25,-18,20,-42,-26,6,10,-21,-2,31,-15,-24,1,35,-58,24,5,-9,-40,11,-5,34,-16,0,38,30,-22,23,21,-9,6,-43),
	(-5,13,18,-6,7,-14,-1,9,0,-2,3,-8,-12,0,-11,-10,-18,-9,8,-1,8,12,-4,8,-7,10,-8,-5,-20,-19,-17,-18,2,5,-11,-11,4,-6,-12,7,4,5,3,13,7,-1,17,-9,16,0,-7,-14,6,-9,-4,8,-11,1,0,-7,-11,15,-11,-1,-4,10,20,9,0,4,13,14,18,-9,0,-17,-15,-16,16,-19,-13,-20,16,-9,12,-4,-2,20,6,-12,19,6,-8,0,-7,-20,0,-12,-2,-16,-11,-7,7,17,-18,-14,14,14,-1,-5,14,-17,17,12,11,6,-9,-20,-4,3,-9,-8,-2,-6,5,-7,-10,9),
	(2,-8,3,11,13,-5,-1,4,-2,-2,1,17,-10,26,-4,-18,17,11,14,-23,-10,-12,-5,0,11,0,-3,16,-3,16,6,-11,-24,23,20,11,-14,-15,-19,-10,-11,19,0,16,-2,19,20,-17,5,-10,13,-21,-15,18,1,-3,9,-20,15,-2,-19,-3,-8,16,-10,7,12,-5,-5,6,3,-14,11,-3,18,-12,-9,5,-21,-24,-14,-19,17,1,17,0,-16,21,-6,19,19,-22,2,21,-6,-13,-10,-25,4,7,-7,-2,8,-11,-5,17,-9,-3,-17,0,-20,-7,0,-13,14,-13,9,1,11,-16,-11,5,-8,15,15,7,3,1),
	(2,-2,-11,-6,-11,-3,4,16,8,3,0,-20,-16,-16,0,6,-6,-4,-14,19,-4,12,8,-22,-8,-7,-11,8,-6,-16,8,-12,-12,11,-4,19,-17,-4,13,15,15,-7,-17,21,-3,15,19,4,6,10,20,5,13,-7,0,-21,-3,23,15,5,21,12,-14,5,0,-5,0,7,23,7,16,16,8,-5,7,20,-20,-14,-8,-1,9,8,13,22,18,-11,-7,17,-17,-2,-15,7,-11,9,-6,9,-9,-6,-10,-13,9,13,8,0,-20,-2,-15,1,14,-10,-12,9,-18,-10,-14,22,14,1,13,-9,-15,-6,12,17,0,-1,-16,-8),
	(-8,-1,-35,26,-25,19,6,44,19,-14,9,-13,24,-4,-17,29,54,-7,-6,19,-2,-18,14,-52,-31,43,11,44,5,-25,-8,-17,13,-18,-20,-14,-11,-7,-6,-22,-29,-28,5,9,-2,14,-15,-1,-6,-5,3,42,-34,-16,22,5,-13,-8,-42,19,-8,25,14,-1,-1,-18,-49,-13,25,-6,19,10,26,22,0,12,-9,8,-5,39,-7,0,43,24,15,-12,-1,-19,-4,-4,4,-27,-31,36,-33,3,63,2,-2,4,3,3,-16,4,-18,34,-12,-5,10,0,3,5,9,-2,46,19,-6,2,-13,13,21,-12,-5,-3,15,-2,28,-2),
	(15,-27,-18,3,4,30,18,38,4,-32,27,28,18,-18,-29,13,44,32,16,1,-20,-38,-23,-3,4,49,-24,0,-1,18,30,-17,38,-2,7,12,0,14,12,0,-19,5,-13,-17,15,7,-6,22,0,-29,12,45,-22,6,11,-2,9,5,-13,-3,17,0,2,-24,-25,-23,14,41,37,-13,9,9,2,34,-2,42,0,6,-29,8,4,5,20,-22,41,-34,-1,7,2,0,-14,2,-14,13,-7,30,19,28,-17,-60,17,5,17,28,-4,42,2,-57,6,-22,-25,15,25,-4,-31,29,3,18,-16,28,9,17,-29,-56,-21,-16,-4,14),
	(9,-52,-3,7,23,33,8,21,29,-43,12,11,8,-23,-45,12,1,6,27,0,-1,-14,-6,-21,-14,27,-9,26,1,19,24,8,-12,-10,3,17,-13,2,43,-4,23,-8,0,-41,-14,13,11,-2,-6,-3,6,-2,10,31,2,-11,-5,-24,2,15,5,3,-25,-35,2,6,2,-15,23,-7,10,20,-6,-10,24,2,16,-10,-38,6,8,-5,-7,1,10,-18,-24,-7,0,22,-3,-12,-23,-25,-19,21,13,7,-34,15,30,1,-29,23,-25,-10,-3,-1,49,-8,18,4,17,5,7,-15,-2,-11,28,3,4,-5,12,-36,-13,4,-4,20),
	(-2,-68,-66,9,29,27,1,13,3,-45,18,-9,42,1,-43,9,-4,44,36,-10,9,64,27,-10,-19,-6,7,2,7,24,15,-9,-23,-19,-4,13,-14,5,48,-30,5,4,-3,-19,-40,6,25,27,-28,6,30,-19,7,32,11,-4,10,-20,12,-4,5,23,9,-8,-41,1,-8,10,21,-22,23,10,-38,-20,22,11,-12,-25,-30,6,-6,-31,25,19,11,-22,-26,-29,-3,5,5,-28,-38,9,-11,25,-21,-13,-32,2,9,-12,-6,32,0,33,-8,8,33,-13,-11,26,-37,15,10,8,-7,27,16,7,23,-4,-28,-29,0,-10,-3,11),
	(-4,-38,-56,36,16,-16,13,14,40,-24,34,-1,26,9,-51,27,-16,28,6,3,32,55,27,4,13,-12,22,1,-9,-6,1,2,0,-23,-15,15,-26,19,28,-28,29,-26,-18,-34,-3,-10,10,-23,-12,-11,14,0,34,12,-7,-10,-20,19,6,-11,-11,-6,-2,18,-64,-25,27,-4,6,17,11,26,-23,-18,17,9,-6,-2,-6,20,-24,-10,-5,4,22,-14,3,-7,-17,-10,0,-3,-27,2,-41,28,5,-25,-75,-22,4,-17,0,13,-3,46,-6,-1,62,-23,10,-1,-16,19,-7,7,-27,2,23,30,15,22,-51,-8,-25,-9,7,-10),
	(-39,-39,-53,28,-2,-16,11,27,37,12,6,-13,31,4,-53,5,-8,42,15,3,-16,59,21,-3,10,23,8,-5,23,3,1,3,15,-23,11,19,7,14,31,-26,8,9,-34,-36,-27,-24,-20,3,-6,-19,21,-1,35,12,13,-13,-12,-12,25,-8,-17,-15,-13,-9,-65,10,11,-2,-17,-5,17,-1,-28,1,19,9,-14,14,9,-6,-18,-30,-10,22,39,-6,2,0,-23,-5,-8,-8,-28,-9,-18,32,-7,-16,-43,3,1,-2,22,18,17,36,17,5,19,-7,13,8,-23,-12,7,-2,-6,16,2,3,12,9,-42,-16,-4,-17,10,2),
	(-26,-56,-41,32,26,13,45,0,4,4,29,-12,18,-12,-48,19,-19,15,5,-10,8,49,31,-3,-4,-6,-1,-14,5,23,1,-18,1,-11,8,-18,16,-14,26,-16,43,-10,-31,-19,-9,-26,-29,-11,-30,7,18,-2,5,32,0,-4,-26,7,12,-4,7,8,-11,4,10,10,5,21,0,-3,8,15,5,-33,-10,40,17,15,22,5,5,-41,-6,-23,36,-22,16,12,-16,-6,4,4,-4,9,-20,35,17,-25,-27,-3,-15,-31,17,17,-13,32,-17,-20,36,0,-17,30,-27,-16,0,38,-7,6,1,16,-13,6,21,-18,-28,-25,-2,-8),
	(-21,-56,-22,14,25,-19,50,-12,16,-3,37,-3,3,-23,-24,33,-26,4,-24,12,-10,-1,7,-8,1,9,8,3,-18,2,8,5,-3,-17,9,15,7,-4,8,-40,20,-6,-34,5,-30,-23,2,4,-24,4,18,12,8,6,19,-16,-21,-10,22,0,10,-23,-6,8,2,22,34,24,-39,18,-3,10,21,-6,-1,38,-5,13,19,-1,-10,-34,-28,-22,23,-17,18,3,-27,2,-2,-7,16,-10,-19,28,11,-23,-27,-4,5,2,3,8,17,4,-6,4,33,6,-4,47,-16,-10,-25,21,-8,36,17,28,19,6,33,4,-18,-3,10,-35),
	(-16,-39,-23,7,17,16,46,-18,21,-16,22,-31,12,14,-15,8,-8,24,-22,13,-39,-19,-8,10,6,26,16,13,1,35,-19,-3,0,27,6,14,-3,-3,-3,-4,15,-1,-43,21,8,7,-12,5,5,-15,5,15,23,13,6,-13,-18,-11,14,-20,10,-1,20,16,31,25,13,48,-12,36,5,-6,-7,-14,-8,28,0,30,25,8,-1,-9,-38,-19,0,-3,0,-4,-2,-16,-28,26,-13,-4,-17,23,34,7,6,27,23,10,7,-6,15,25,-26,-10,13,14,2,28,36,1,-4,28,-3,14,29,7,6,30,-13,-11,-26,33,13,-1),
	(1,-7,-3,17,-1,-2,8,-20,15,4,25,-10,-36,-30,-21,47,-5,9,23,-2,-9,-50,24,30,4,15,-4,-13,-9,10,1,-6,10,-8,8,18,16,-22,1,-6,18,-7,-19,-17,42,0,5,-21,22,-3,-4,33,8,10,15,-18,2,9,-8,-9,15,-10,14,20,-19,27,36,23,6,35,5,-18,-28,2,11,37,11,25,2,34,3,-3,-6,-8,22,-14,18,-8,-22,-29,5,1,-6,1,-20,23,12,-22,1,22,-12,-5,44,13,16,18,-23,-11,12,-9,-21,53,14,13,-17,3,34,7,5,-1,3,13,-5,-19,-29,10,18,-12),
	(-6,5,23,12,-12,17,7,-1,-5,18,-17,-21,-21,-17,14,41,-14,17,13,-15,4,-23,-10,4,-6,-1,13,2,-37,50,-18,-24,2,-1,-8,11,20,-1,-38,-11,4,1,-19,11,20,-12,13,-23,-9,19,-9,-14,-8,0,10,3,-24,10,28,-3,2,-27,-4,-6,-29,14,45,30,8,25,9,-3,11,-20,-23,13,29,17,-5,-7,-20,22,-33,4,-20,-18,1,0,18,-2,-18,21,6,4,8,25,-14,-5,-6,28,-7,17,30,24,23,17,-7,7,-24,12,-8,36,16,-9,-15,13,6,40,13,28,21,-16,-15,8,-14,27,39,-4),
	(20,7,-8,21,16,22,-15,-7,0,8,-10,1,-24,-40,-1,13,6,28,-2,14,-1,-29,-5,20,-8,7,-4,17,-3,3,0,-8,0,20,15,21,-18,-26,-26,-2,18,2,24,3,18,0,-4,3,5,-11,-3,-2,-17,-21,-16,-31,-21,-6,-14,6,32,-16,0,3,-18,28,47,36,-33,-9,5,-11,-17,15,8,-1,-12,14,-17,1,-1,24,-24,15,25,-9,31,4,0,6,-6,24,-10,24,6,0,-5,1,-1,-1,-22,0,23,21,29,0,-6,8,-26,-1,-13,28,31,-11,-12,24,23,25,-23,13,16,-27,12,23,-57,33,21,-6),
	(33,3,20,2,-6,-5,-36,-15,-2,5,27,12,-11,-30,-3,22,-1,17,16,6,23,-29,16,10,-6,-6,-4,14,1,33,-33,2,26,36,10,-4,22,16,-33,10,5,-3,14,11,-1,-2,2,-15,-5,-8,-38,18,-22,14,0,-20,7,23,7,-16,15,6,-24,10,2,24,18,26,3,-11,7,7,-29,6,3,4,-14,3,6,-16,20,22,-34,17,8,-37,33,-21,20,-20,24,8,2,19,22,-7,16,-15,-15,-14,-31,16,38,13,1,22,12,-14,-29,16,19,33,4,0,-2,5,17,27,3,9,13,-8,17,13,-56,12,2,1),
	(5,6,-7,-4,-8,-14,-41,-15,-21,8,8,14,-10,-41,-10,-6,19,-13,14,23,0,13,36,-16,17,5,9,5,-9,39,-26,-4,-6,33,3,29,-2,-18,9,-4,10,17,20,22,0,-5,-15,-25,19,-4,-33,16,2,-21,-11,-7,19,19,12,-13,18,7,-17,-23,-13,2,-17,10,-10,8,19,8,-13,11,18,-28,9,2,-7,14,0,15,-43,-2,12,-16,19,-12,20,15,9,36,21,5,-13,-25,12,6,20,-37,-3,2,20,-7,13,-3,-5,0,9,-14,-6,12,13,-3,13,3,0,14,-12,15,26,-32,2,48,-39,40,9,-8),
	(27,26,-16,4,-5,3,-25,11,2,-7,19,41,-7,-36,24,20,-15,13,-17,-15,-8,30,10,-32,7,15,15,9,13,37,5,-13,19,20,-4,0,13,0,13,7,17,22,-11,1,17,-6,0,-33,5,12,-11,11,-23,13,-12,-21,17,14,2,16,13,24,-28,-7,-3,10,-33,17,19,-17,19,9,-41,-7,9,-24,4,7,-4,8,0,27,-53,19,16,3,16,-14,44,20,12,0,37,-5,13,-34,16,-18,11,-19,-18,13,20,8,-24,2,2,-14,19,5,-11,47,14,15,-7,0,2,-12,-12,22,14,6,-21,35,-42,17,8,-12),
	(24,47,7,14,-3,11,-17,-13,-11,8,40,36,-12,-21,-18,27,4,20,-2,4,16,35,28,-13,3,-6,8,-2,-14,8,16,-5,-13,-2,-23,16,4,19,24,0,9,17,-15,0,31,-6,-33,-16,8,9,-22,16,-1,0,10,2,16,4,-29,-8,-17,18,-18,-16,-12,2,-71,0,-7,-17,25,7,-5,-15,24,-45,-12,-5,-15,-4,12,4,-41,-24,24,-24,-11,10,19,13,-2,16,34,-3,-13,-38,13,0,-14,-27,-15,-5,0,28,-19,-2,-4,-35,-14,-15,-2,4,20,6,-12,5,25,25,15,18,16,-28,14,14,-46,9,27,7),
	(6,26,-15,28,2,22,-19,6,12,4,48,30,8,-30,-27,33,3,17,14,13,-17,36,-1,-18,-4,20,27,12,-4,14,31,-30,2,-5,15,-1,-33,-9,23,21,27,-12,8,2,24,-8,-4,-8,0,-34,-29,-8,-10,-8,-3,-2,-11,12,-10,-8,-31,22,-21,11,18,2,-78,0,7,14,2,33,-2,-4,14,-28,-12,10,3,-27,25,0,-48,-49,13,-24,-6,0,24,27,12,5,6,-17,1,-52,-13,-13,-14,0,10,1,-12,30,-21,-6,11,-8,6,-30,13,28,0,7,-19,-8,-9,10,-32,-6,20,-23,8,10,-37,10,29,12),
	(2,46,-31,0,10,30,-15,29,-15,9,21,54,-20,-40,0,23,24,4,-1,19,-29,13,4,-43,-27,20,3,6,12,-7,-9,-31,-9,6,25,31,-26,27,0,34,0,-24,-14,-5,0,-8,-16,24,1,-21,-23,-1,-32,6,-1,-24,-36,-1,-12,0,-29,11,16,8,-16,-12,-89,17,-13,0,0,16,-51,1,45,-38,9,16,-32,8,-19,-7,-30,-37,13,-3,-15,0,-2,18,25,-27,-22,-36,-36,-50,-20,-21,-45,-2,-2,15,-51,24,8,-28,-6,-38,-9,-29,3,8,17,-8,-20,-10,-20,12,-22,30,23,14,-9,10,-7,13,21,-6),
	(13,22,8,-3,34,33,-38,5,-11,7,19,44,6,14,-17,-4,17,-15,-35,-12,0,-15,24,-27,-27,27,27,30,-6,4,23,-4,-41,-4,6,7,-10,8,11,-17,16,13,9,22,31,-10,-37,20,-11,-27,1,15,-46,45,12,8,-39,-18,-8,13,-41,18,6,-5,-19,-34,-58,-29,-14,-27,10,0,-77,-12,25,-31,-11,-8,-1,-26,-8,-4,-10,-20,35,1,-36,27,4,1,18,-11,1,-5,-1,-17,14,-32,-37,11,-6,-6,-52,-2,-22,-14,3,-34,14,-39,0,12,11,16,-38,-31,-3,1,-49,19,-8,-2,11,2,-44,6,-5,13),
	(40,7,1,5,59,52,7,10,11,14,19,5,2,9,-52,9,19,-1,-21,-8,-15,-21,24,-21,-43,8,16,11,18,4,16,-47,1,-11,-8,8,-10,13,-33,-14,16,-4,3,21,43,-33,-29,7,-9,-31,-43,3,-42,26,-18,30,-61,-16,-26,-5,-37,7,4,14,11,-4,-31,-4,-14,-21,19,-25,-50,8,-2,-4,-1,-21,-24,-4,-8,14,17,6,2,11,-37,-2,-21,-37,-5,-47,3,-27,-4,-43,-24,-2,-71,23,11,-6,-76,6,-18,0,19,-42,-6,-12,-6,21,5,10,18,-46,-33,9,-45,-17,-5,-14,4,21,-14,6,-5,-4),
	(-16,18,14,28,30,27,-6,19,0,4,37,8,-3,35,-36,1,12,14,-20,14,-27,-54,31,-8,-7,19,2,22,-16,-14,10,-26,9,-9,-22,-16,1,8,-19,-7,-7,-5,-16,-3,19,-15,-18,0,-20,4,9,35,-20,12,11,9,-19,-15,-8,5,-58,0,37,25,-34,-23,-4,-15,-8,-16,13,-16,-28,3,0,7,-11,14,-21,-1,-20,42,25,-21,0,-12,-6,6,9,-32,-36,-5,-17,8,-4,-31,25,0,2,-3,16,0,-48,27,0,-8,-4,-42,-30,-26,18,25,-15,-9,16,-10,-39,-5,-44,0,15,-14,-12,-9,-43,-17,-9,22),
	(38,22,24,-1,-11,-2,-16,12,-3,6,17,-15,45,30,-5,0,-1,12,-33,3,8,-29,2,14,10,16,13,35,-32,14,41,-45,23,-1,-3,-23,-15,16,1,1,20,-15,1,7,58,-38,-40,-31,-19,-26,-11,48,-20,48,2,40,-12,2,-25,4,-44,26,-10,0,26,-11,-23,-17,-8,-19,23,24,-8,-15,-5,-5,45,-9,4,-17,-19,26,0,-16,37,6,17,12,-18,-47,-43,-18,1,-37,15,1,9,34,15,12,0,0,-40,1,-19,-7,-4,-52,-51,-14,-1,18,1,-21,27,-34,-45,2,-10,22,33,20,16,21,-36,-18,4,-28),
	(23,9,52,31,23,-11,-4,3,-31,-43,35,-22,58,30,23,15,-26,29,-9,-9,17,18,1,14,-2,16,-3,35,-2,-17,69,-34,-2,-10,1,-38,18,20,-23,8,-2,-31,-8,11,5,-13,-69,-3,-27,-52,-51,14,-34,25,56,41,-4,-16,-2,12,-22,26,27,-27,28,11,-5,-53,-4,-24,-15,-15,-35,-3,20,-11,50,32,11,-21,-14,15,0,-16,7,13,0,8,-39,-37,-27,-8,-11,-27,2,4,-15,-3,-2,-5,41,-32,-16,-1,10,-16,-11,-45,-49,3,-3,45,-65,-46,-14,-17,-47,-41,14,-27,26,18,23,14,-18,-8,12,-23),
	(0,-2,21,1,6,-1,8,-10,7,-29,7,-18,-7,29,15,2,-7,9,-7,-10,7,30,-12,8,-4,12,1,-25,-6,10,38,-6,-17,-6,20,13,24,14,-7,-14,-11,-11,-9,-15,-9,-1,-2,-4,-19,-39,-27,10,18,24,45,0,-10,-18,12,-5,-17,20,-26,1,25,-5,-36,-23,29,3,8,-7,-24,-4,-17,-17,-3,12,-11,-21,16,13,-31,39,18,19,-26,-23,-10,1,3,-25,-11,-29,8,-23,-23,-27,-39,-4,-4,-19,-16,-9,12,-28,1,-17,-2,11,20,4,-51,-30,1,-26,-15,-46,-19,-38,17,-3,-17,49,-24,5,0,-13),
	(-11,39,-1,-7,44,-8,-36,6,-23,44,-13,31,-26,31,-13,-11,-19,-12,-19,-11,-16,-17,6,5,31,-18,18,-32,23,16,14,-18,-20,2,19,24,15,35,14,5,-20,29,-14,-14,-8,33,-17,26,6,-53,6,22,4,28,-17,-37,-17,-11,-20,-11,7,-2,-20,4,45,10,0,1,23,1,-28,27,29,-23,0,-11,-14,-4,-35,-18,8,3,-3,44,1,34,29,44,-37,43,25,-16,36,-21,-48,-28,0,-35,26,-13,-21,26,-33,9,0,-37,-18,-9,15,-19,-28,7,3,-16,-24,-26,-21,41,9,-7,18,16,-26,-4,-29,22,-22,-24),
	(6,-12,5,4,-7,-6,-11,4,-14,16,12,3,-20,0,-19,11,-16,6,-14,1,-13,-19,-16,6,-19,17,-20,8,18,-1,-12,9,-18,10,-9,14,-10,17,14,10,12,11,14,-7,-7,18,-4,-14,6,12,-18,8,-6,-20,4,7,1,15,20,13,2,21,-6,4,17,-1,-16,-3,19,3,-6,7,0,7,3,-4,-15,17,-20,19,11,-4,7,2,-9,-18,-16,-9,-12,-19,-11,11,-8,-16,20,17,-19,-12,10,-2,19,-21,6,-19,-5,20,14,18,0,1,-17,20,-20,-16,18,-9,-6,14,3,4,-11,-7,-8,-14,12,-14,10,-11),
	(9,9,13,3,-18,13,-10,12,5,19,-18,-19,-5,16,-2,15,15,18,-8,16,19,-15,14,-1,5,1,-15,-18,15,8,20,4,-15,-3,1,9,-18,-16,20,11,-3,-18,-12,16,-12,11,0,2,13,10,-7,-19,-14,9,-9,-3,1,9,4,-5,-1,-18,-8,-12,14,17,-14,1,4,-13,3,-14,-20,-4,-13,6,-1,0,10,10,-12,19,-2,7,-5,0,-8,6,10,-18,7,12,16,15,-16,-18,-2,-14,20,6,14,-7,-1,10,-17,4,-8,-18,-6,3,-19,10,-1,15,5,1,15,1,-15,16,6,-9,-5,16,3,11,-14,1),
	(19,11,3,-10,7,1,7,6,18,-17,7,-12,17,11,7,17,-11,11,0,20,18,-6,-4,0,12,-5,14,-14,0,-14,15,-17,-20,13,12,17,-18,-6,2,-4,-19,-9,12,-18,-12,16,-11,-3,0,0,5,14,11,-8,-8,-20,20,-4,-13,-7,5,5,-10,-11,10,14,-18,14,-6,-16,4,0,-17,10,14,17,-5,-16,18,6,-18,-2,6,18,18,5,-4,10,16,10,7,-11,-8,-5,-16,15,-9,17,-11,10,-9,19,-4,-8,-5,18,6,-14,-9,-16,11,2,-9,-7,-9,10,-16,16,-9,-19,20,-7,-18,7,7,14,0,14),
	(-4,-10,-23,22,-15,10,-32,36,21,-14,32,22,-12,-36,-20,7,20,7,-10,22,-5,-12,2,-27,-6,14,-3,-11,48,22,-17,43,9,-3,-18,31,-12,36,-1,16,-27,-17,-9,-10,-2,-13,6,1,13,32,27,6,-32,0,39,-33,-45,16,-34,18,31,55,17,-2,-23,-8,-34,16,29,-28,14,31,26,-5,30,8,-26,4,-33,47,-9,22,-16,4,12,-13,-27,12,2,6,-2,9,-33,-26,-42,-10,34,-8,8,-10,21,0,1,33,-8,15,-11,-14,14,-18,-41,-16,21,19,58,8,12,8,-3,26,-5,-22,-12,-25,-2,-11,-2,-13),
	(16,-19,-4,4,-21,18,-11,20,-4,4,-2,43,-14,-6,-36,29,43,-32,-11,9,-31,-25,-24,-28,-28,43,-32,9,14,26,25,18,57,-14,-13,30,2,2,15,8,9,-6,-26,-29,47,-10,1,-11,21,23,17,33,-36,20,23,-35,-11,11,-51,-8,19,-3,-13,-12,-39,-35,-2,42,47,2,36,24,10,-7,17,33,-6,21,-51,-5,-29,36,15,-13,42,-55,31,40,3,41,27,0,-15,-40,-19,9,75,26,-17,-29,-12,7,17,24,-7,-3,-10,-27,3,-25,-18,-3,34,41,9,2,54,4,-5,32,26,8,-47,-9,-54,-14,14,-3),
	(12,-73,-19,6,-29,22,-33,11,30,-28,1,11,-11,-26,-27,18,18,6,30,16,21,17,-42,-29,6,16,-7,-8,-9,23,38,32,-3,-6,32,-13,9,32,8,12,13,15,-11,-57,0,-9,3,-20,19,20,1,5,23,33,-2,-18,-28,-2,-44,17,11,-5,-42,-30,-54,-1,11,14,48,-2,-3,30,-21,-2,10,33,10,-7,-24,7,-42,12,-35,26,12,-19,39,45,19,29,7,-30,-5,-54,7,-16,28,6,-33,-4,-4,8,-28,-5,-18,7,0,-15,12,-29,-16,-24,17,2,37,-24,4,1,6,5,24,0,-27,7,-45,-4,4,2),
	(-1,-62,-12,5,-23,-8,-18,-10,4,2,-16,11,10,21,-38,-9,3,21,13,-4,10,74,2,-34,-9,-1,-34,-4,14,9,21,29,10,-18,22,3,20,20,35,5,13,46,5,-38,-23,-13,-27,9,21,10,8,10,-4,1,13,-18,-22,17,-20,18,18,25,-28,-28,-52,0,-16,36,16,12,0,25,-14,-10,16,28,15,-18,-1,-10,-1,-15,0,25,9,-28,7,26,-13,-13,4,0,-47,-37,-7,12,-26,-14,-20,-5,-16,-8,-19,-6,-5,-14,-19,12,24,-28,-15,-8,-9,8,-22,-8,-15,0,7,14,42,-4,-43,-34,-16,-23,3,-5),
	(-20,-34,-3,-2,-7,-3,11,-3,-8,-1,20,-4,14,44,-53,21,5,-1,3,41,2,49,43,8,-21,-29,-4,-12,-1,14,-32,21,-9,-35,20,10,2,8,31,-16,-15,-2,-28,-75,-31,-1,11,-15,-2,-4,24,12,3,18,0,-7,-38,36,-5,6,11,18,3,-14,-83,-20,10,9,56,18,2,22,-40,-12,-15,54,7,12,8,-2,-1,-24,8,13,24,-9,17,1,-9,2,4,4,-36,-8,-23,30,-36,-1,-51,-2,-34,-6,-19,-8,-5,12,-17,6,27,-2,8,0,-39,5,12,10,-22,9,5,29,39,-3,-46,11,-16,-5,18,-14),
	(-22,-41,-20,20,-21,-22,8,7,32,1,9,-6,29,19,-37,14,15,6,-4,6,10,53,13,8,0,-5,-20,0,25,-3,-23,7,-8,-33,-23,1,9,-6,46,-2,5,-8,-38,-37,-25,14,-22,-39,11,-9,15,-4,0,11,-1,22,-32,8,44,-17,0,3,24,18,-37,12,14,4,29,6,11,21,-66,-19,-13,33,-20,28,29,13,-9,-1,37,12,28,36,35,-19,-15,24,5,-7,-25,-15,-33,19,10,-12,-26,33,-40,-19,4,17,-4,-3,-15,-14,40,11,12,21,-33,-6,-4,7,-20,15,3,34,1,-10,-5,-1,-2,-44,16,4),
	(-8,-70,-16,13,-14,-9,40,14,0,-5,8,-7,-8,-1,-49,21,14,20,10,5,6,43,-1,20,-10,27,14,-3,13,7,-15,-6,11,-41,-27,20,0,-22,28,-24,1,3,-45,-21,2,-11,-15,3,-6,-15,20,37,-3,-6,-4,-1,-39,-5,2,0,-35,-26,7,5,17,18,23,-3,-6,-1,-10,-4,-24,-35,-19,54,8,33,-9,29,0,28,2,-13,12,8,7,3,-15,6,-21,34,24,-15,-34,21,18,9,-26,13,-42,-20,3,16,9,27,22,0,25,-12,19,23,-7,-14,-8,5,16,7,21,17,1,26,-14,22,-10,-34,-3,-8),
	(-35,-94,-19,4,25,-10,17,-1,3,5,23,-11,-14,4,-38,33,-20,19,1,20,21,18,6,20,1,-13,28,25,0,36,-6,-25,23,-33,-14,1,-11,14,23,-10,12,20,-29,0,16,6,0,-18,0,-29,40,5,1,-18,5,2,-20,24,10,-10,-23,-17,-8,18,0,-3,32,17,9,23,-13,15,-22,4,-19,30,14,24,-18,-2,6,9,-36,0,16,0,2,4,-14,15,0,10,2,5,-42,11,20,-9,6,-19,-35,-29,14,40,12,13,1,-11,20,21,3,2,-10,-26,-8,19,2,37,-9,-9,-5,19,13,4,-13,-28,0,-39),
	(-4,-47,26,14,6,-12,30,21,8,16,14,-4,-16,17,-10,9,1,10,0,4,-10,-5,26,9,31,2,34,26,-16,49,-5,-15,15,0,0,17,-4,10,14,25,28,-13,-32,-9,0,4,4,-31,23,-22,5,22,-2,24,7,-14,-11,-1,17,-17,-2,-8,28,9,27,0,15,-1,6,11,-2,-5,-18,10,-5,54,-9,-5,8,34,7,-5,-47,6,23,-2,33,22,0,7,-21,24,3,7,-36,43,27,-25,26,21,-13,0,-1,7,5,1,-12,-31,10,5,11,38,22,-3,-16,28,-2,26,38,37,8,12,12,-18,-7,-27,32,-1),
	(-10,-52,5,9,-7,-24,3,1,15,4,26,-12,-24,-24,-2,43,-11,11,6,15,8,-25,15,10,12,-23,20,33,-13,19,-9,-14,13,-14,-23,18,-11,-4,0,-9,14,-5,4,-5,31,2,24,-59,-5,-2,-5,48,20,22,2,11,1,6,19,17,6,3,38,27,13,11,11,23,-9,4,-5,17,-18,20,-26,25,6,9,6,25,-12,0,-17,18,36,-13,30,4,-8,16,-10,5,-28,-1,-25,3,9,10,20,26,-4,-12,38,30,17,22,9,-12,-17,-12,-12,20,18,-7,-23,-3,5,48,38,47,20,31,-13,-22,16,-24,5,22),
	(0,-33,-6,13,3,-15,36,-16,-20,6,39,2,-9,-19,-13,24,18,20,11,10,18,-37,0,52,18,17,17,24,-13,49,2,-12,0,23,-16,-4,-22,-21,-11,-17,7,31,5,25,10,15,7,-14,2,-9,0,5,11,7,5,10,-11,7,9,-8,-8,-13,11,2,8,-4,1,15,6,1,6,-13,-24,-9,-29,20,15,-5,-3,16,26,2,-19,14,37,-19,27,9,-10,12,-23,29,-3,24,-16,5,23,-32,-2,-4,-10,17,37,9,9,15,18,-16,-37,-13,8,50,0,9,-37,-1,3,12,12,18,0,22,17,13,-23,-7,13,-8),
	(-18,-8,-1,16,12,-19,11,-15,-10,19,27,19,1,-26,-18,15,7,13,20,-4,31,-15,8,8,-1,-15,31,19,15,28,-26,-35,-2,28,5,0,-1,-4,-13,-7,-2,-2,16,26,5,-8,24,-40,7,-9,-28,37,6,-19,-13,-20,21,26,-12,-7,0,22,4,21,-3,18,-11,-2,-16,10,0,-10,-33,-3,0,4,8,-8,3,-1,-6,0,-19,21,22,-36,21,-28,12,4,0,40,-14,7,0,-12,-3,0,-10,-29,-23,28,22,28,24,28,-2,-13,-2,5,23,7,12,26,19,10,0,3,29,13,13,-16,1,-17,-22,0,28,9),
	(16,19,18,13,12,4,-11,-31,-9,16,10,51,4,-31,12,7,-13,-4,4,-11,1,-26,0,3,5,-16,22,6,-5,39,-20,-2,10,20,-12,2,-4,0,-11,-3,-8,11,17,5,29,8,9,-26,22,-8,-26,13,5,-15,13,-12,22,10,-2,-18,-14,9,-18,20,-17,24,-17,-7,-7,23,-16,17,-23,4,-5,1,-19,-3,-11,21,-1,28,-21,-3,24,-3,27,-22,9,-19,22,36,0,-2,2,-25,1,12,-9,-38,-40,22,26,18,-4,3,18,-7,-5,-6,8,35,26,11,15,1,15,17,10,29,12,-11,16,2,-31,25,24,23),
	(6,45,-22,2,28,-12,-38,0,-15,0,4,59,-9,-14,-1,4,-22,-2,17,-15,33,18,0,16,-2,4,30,-5,10,36,-29,-5,10,12,-11,16,-22,-4,-9,16,23,24,31,25,2,-37,5,-8,13,11,-4,-4,14,-8,-15,-19,11,7,-5,2,13,-13,-18,-4,8,7,-46,0,-3,13,3,24,-15,-8,-13,-14,-14,20,9,8,30,25,-32,-18,44,-16,29,4,10,-9,26,27,7,9,12,-3,-4,-13,9,-27,-20,22,-12,28,-5,-14,-3,-7,12,-12,-2,18,13,30,3,12,-2,17,-13,-1,15,5,4,19,-35,23,14,-5),
	(23,31,5,26,2,2,-10,-3,-2,-3,48,42,-1,-32,-8,26,-23,8,-5,11,22,18,19,-3,-2,9,24,19,5,-4,-8,-22,-13,4,-5,19,-17,3,32,16,-9,19,-8,9,13,-24,26,-25,23,-4,-24,16,-6,9,-18,0,11,-15,-12,-13,-30,-11,-24,-6,-7,14,-77,4,-13,-1,-4,11,-20,3,0,-11,16,11,-24,0,4,11,-41,-4,32,-23,22,7,22,-22,22,23,15,-2,7,-25,7,8,-44,-23,-49,33,-27,12,4,20,0,-11,3,-6,-7,10,15,-5,8,5,-1,2,7,1,2,-10,1,10,-12,13,27,9),
	(14,46,-14,6,21,14,-22,26,-9,-3,29,50,-14,-45,11,13,-26,-7,-6,-9,23,44,-12,-37,5,4,27,-13,-2,16,18,-12,-14,9,-23,20,-24,-3,19,-16,25,-17,-1,41,30,4,-18,-20,-10,-6,-33,8,-29,-1,-19,15,-8,4,-2,-8,-19,0,-27,10,50,-1,-75,-6,-17,-1,20,28,-31,11,5,-30,-18,30,-1,-19,7,6,-54,-29,17,-24,18,-18,2,-22,13,11,-3,0,15,-54,-2,-1,-44,-17,-27,-9,-11,32,-19,24,4,0,-9,13,16,11,13,20,20,-18,4,0,17,12,13,-11,-14,39,-47,24,5,30),
	(0,45,-28,1,37,34,-22,21,-10,3,27,31,-11,-38,-15,21,4,7,-2,-16,-5,48,14,-25,-20,62,-11,-5,-15,0,-9,-34,4,-4,11,30,-13,9,13,20,-4,-17,14,33,58,-8,-14,-22,11,10,-18,6,-33,13,-20,4,-22,-6,-23,2,-34,16,-30,14,35,-28,-89,33,-19,-26,26,3,-25,-1,45,-22,-3,21,4,4,7,26,-34,-23,6,-21,-2,4,53,-9,-13,9,-26,-23,-4,-21,-4,40,-45,-19,0,-10,-50,8,-23,10,0,-35,0,-1,0,15,50,9,-16,-17,12,-4,-29,-4,3,-5,0,32,-72,21,-3,34),
	(17,16,7,0,31,48,-28,25,2,19,51,-5,-6,-34,0,21,2,-13,7,1,-33,45,11,-51,-14,41,13,19,-5,-21,26,-7,-25,-3,10,8,-26,2,10,0,-9,-32,11,19,45,-8,6,5,-16,-27,0,-4,-28,9,0,14,-40,4,-33,17,-47,-13,6,12,-11,-21,-79,8,-29,-13,29,-3,-71,-27,40,-31,32,4,4,-6,17,13,-46,-67,-2,-18,6,5,20,-7,-3,5,-19,-19,-11,-29,-5,18,-14,-30,-2,4,-38,2,-2,-6,-4,-31,30,-5,22,5,13,0,-34,-12,-10,-6,-21,-12,-7,1,-5,37,-52,8,12,9),
	(-6,19,5,8,29,26,-9,22,4,21,27,-13,-11,-22,0,5,-12,0,4,-7,-24,15,-11,-42,-20,22,-16,26,-13,-2,8,-28,11,-16,8,14,-22,0,-10,-27,1,-22,0,44,21,-29,0,3,-15,-9,-41,10,-28,27,-17,16,-54,3,-36,19,-49,0,-22,1,-44,-7,-51,-9,-17,-24,36,3,-29,-33,47,-32,6,25,12,-21,6,30,-14,-14,-2,1,-5,5,-11,-20,-15,-34,0,-43,-16,-33,-5,0,-24,-12,8,-4,-40,18,-15,1,24,-12,-23,-40,6,23,29,-11,-13,-32,13,-32,-35,22,-1,-4,-15,29,-16,0,-16,27),
	(-3,20,-13,-2,35,51,-5,19,26,-7,31,-14,20,18,0,21,11,3,-14,-20,-55,-49,39,-11,-13,49,15,41,-24,-11,5,-51,8,-3,-10,-7,-7,15,-4,-23,-1,-52,3,45,39,-26,-27,-2,-17,-38,-35,30,-35,13,5,34,-27,-35,-33,9,-44,35,16,16,-12,-26,-29,-10,-47,-3,13,-26,-45,-16,-8,-21,17,-5,-4,2,0,48,-26,-3,-18,24,-21,-19,2,-37,16,-33,-12,-2,20,-20,8,35,-28,3,-5,1,-47,-5,-26,-9,8,-29,-37,-42,3,38,2,-41,-6,-23,-2,-20,-31,6,10,-13,-7,4,-10,-5,0,12),
	(-5,7,-9,36,-44,19,-8,50,10,-28,31,-12,25,34,-13,26,-30,49,-23,0,15,-13,1,-22,-5,40,18,32,2,-32,46,0,20,-20,-25,-2,-12,-12,-26,-47,-29,-47,0,14,33,-26,-15,8,-32,-6,-27,33,-13,26,-8,22,-49,-12,-7,6,-47,20,23,3,4,0,-40,-19,-33,-5,22,-21,-12,-10,-29,-6,26,3,-18,-9,-33,48,-1,-17,10,-30,-9,-3,-2,-50,-26,-3,18,-12,44,-20,-14,30,-31,4,38,23,-29,18,-36,22,25,-5,-38,-19,10,13,6,-19,14,-11,0,3,-5,-2,23,8,3,17,-29,-8,14,-1),
	(46,25,23,17,-51,8,-10,57,-17,-41,39,-4,42,47,0,24,-18,36,-26,11,14,-32,-23,10,30,26,1,40,-14,-29,61,-19,58,-4,-9,-41,-1,7,-27,-32,-9,-31,-1,9,64,-27,-33,-25,-30,-5,-35,25,-32,46,12,21,-26,-31,-15,-14,-41,23,0,-12,9,-1,-29,-2,-26,-28,10,0,-12,5,4,40,57,16,-25,-15,2,50,-15,-55,19,-21,6,19,-14,-30,-27,11,18,-33,22,-19,2,42,2,4,24,-6,7,8,5,-7,13,-47,-8,-21,15,11,19,-53,4,-40,-7,-16,-13,-9,29,8,22,29,-41,24,18,-10),
	(24,15,21,23,-41,-22,-10,3,-10,-32,-2,8,48,39,5,-6,-12,17,7,-5,8,25,-27,-10,19,5,-19,22,-23,7,80,18,44,4,-11,-17,19,19,-12,-3,-16,-17,-26,-7,37,-27,-56,-38,-2,-21,-71,-7,-32,68,29,8,7,8,-6,3,9,9,-10,-6,27,6,-58,2,8,0,33,10,-17,-2,19,20,44,26,-11,-27,17,42,-31,-13,-1,12,-3,-2,-20,16,-21,12,-18,-59,25,-6,13,63,-4,8,-1,-29,-2,1,1,-33,-16,-32,-3,-27,-1,42,-7,-1,-25,-33,15,-34,17,-5,20,18,-16,-14,-48,7,-14,2),
	(8,8,30,14,-9,1,7,29,9,4,38,20,-10,50,5,24,-36,-12,-6,-19,-9,14,-32,-1,4,8,-5,-25,0,-13,24,-24,5,-27,-13,0,0,3,-20,12,-22,-29,1,-10,15,0,-37,16,-13,-22,-21,27,12,39,27,10,3,-2,-6,-11,-26,-12,0,-18,5,22,-8,10,11,-21,-28,6,-15,-22,0,13,22,-5,-30,-15,8,24,-33,25,22,-7,-11,5,-21,-4,-22,3,19,-46,-31,-21,-6,-17,5,-9,-1,11,-12,-18,-1,-18,-19,-3,9,-3,-6,-11,-6,-16,-16,-11,-11,-8,-15,-8,48,18,-10,-6,-36,24,22,5),
	(1,38,14,0,39,-16,-38,-27,-22,5,8,5,-3,38,-30,-21,10,-23,1,-1,14,-16,-27,-9,-6,-2,19,-11,4,11,5,24,-19,3,13,7,2,16,20,17,-2,32,-35,13,-11,16,-32,52,-8,-41,-16,-5,-4,-3,16,-29,-11,-33,-28,11,-7,-5,-31,-13,21,4,-26,-21,17,-5,-23,5,23,-17,-8,17,1,-39,-35,-29,2,-4,0,26,30,18,9,36,-10,13,15,-34,0,-5,-41,-21,17,-31,45,-7,-30,13,-33,-28,7,-47,-26,-45,28,-16,-24,-22,-35,-14,-15,1,-38,35,12,28,37,34,2,5,17,8,-37,22),
	(-18,0,-20,8,-20,16,0,6,-16,-4,-10,9,10,-10,1,-9,18,3,0,5,18,-20,0,-2,15,-6,16,3,20,-13,-8,18,3,-11,-18,13,-8,17,-1,-8,-14,-14,0,0,-8,15,19,-2,3,16,1,19,-20,9,14,-14,15,-10,0,-4,16,7,-5,-16,-2,-2,5,-13,0,-19,-19,-12,11,18,-7,-5,-10,-3,0,14,10,-2,15,17,10,-16,5,-2,-17,11,4,-15,0,-10,-5,-13,-15,-4,-19,1,17,10,16,-19,5,14,12,5,9,7,1,-13,6,-14,-18,-13,-9,4,-5,14,17,10,3,-2,-2,0,7,19),
	(-6,-8,8,-6,18,-5,9,13,16,14,3,4,0,-2,7,-10,9,19,3,-20,-6,-14,-4,14,-12,6,-6,5,4,-11,-10,-9,17,19,-2,-3,15,-17,14,-18,19,7,19,-16,11,0,-4,-8,0,3,4,2,-11,0,-17,-15,-2,16,0,18,3,5,-6,16,9,-6,17,2,2,20,-5,-6,1,-9,6,4,14,-18,19,15,-14,-19,-8,-8,20,-11,2,-15,18,2,18,-1,-11,4,-9,12,-10,14,-3,6,16,-20,13,15,7,-7,-16,-16,-12,-20,-4,-1,-6,5,5,7,-19,3,20,1,-10,16,10,-20,3,3,9,12),
	(2,-3,18,-5,-18,16,0,3,10,11,-19,20,-5,-1,19,6,-16,-15,-20,-5,-14,-13,-13,1,-5,-5,-11,13,-2,3,-6,-18,6,8,4,4,-16,-1,6,-1,5,18,1,13,-11,-9,15,11,-15,-7,7,-2,-6,11,20,10,14,-19,11,-10,-5,-3,14,-18,-14,20,11,-8,-7,-5,-1,10,3,11,-14,8,13,-16,-1,-11,-17,-14,9,-18,3,5,-9,9,-14,-19,0,13,18,-2,-4,-1,5,15,2,1,-3,-2,-20,11,14,-14,0,0,-11,16,14,-12,13,-15,-20,-12,-1,4,-19,-16,-17,5,-19,-1,-18,1,-2,3),
	(-10,7,-1,-18,17,0,-22,29,7,8,17,1,-12,0,-8,-18,-1,-7,24,-4,-25,-1,8,-42,5,10,1,6,42,20,-33,39,18,2,4,34,-7,25,33,54,31,-24,-8,-32,-8,17,10,-14,23,32,31,19,-11,28,19,10,15,2,-14,-2,8,3,14,14,-18,-15,-40,-7,8,-9,13,41,29,2,-3,-11,-10,-11,-24,0,-15,5,17,31,-9,0,-19,22,-3,4,-16,25,34,-9,-26,20,-14,-27,7,10,-17,-22,6,7,4,-18,-21,9,18,4,0,-18,7,16,50,-7,10,3,-2,-6,-11,-43,-12,13,-26,-3,0,19),
	(-10,15,-3,-43,-30,-51,-29,29,-31,-15,-42,52,-58,-3,4,-12,50,-47,17,20,-31,-9,-10,-26,-18,-26,-12,-6,1,22,-17,26,44,21,-39,-8,0,21,39,63,25,-41,-25,-30,30,5,-6,-33,58,16,0,-3,-8,40,35,-47,32,21,0,-9,22,29,-19,-16,-8,4,-35,4,48,8,10,46,22,-7,37,-2,-5,16,-41,23,-4,0,-12,47,10,5,9,47,13,17,-23,1,10,-29,-16,13,28,3,31,6,-15,23,1,2,-44,-12,-3,15,39,-33,0,-16,15,39,13,2,34,46,-31,23,-6,-31,-21,-14,-31,6,-11,22),
	(-37,-25,1,-45,-16,-35,-9,-10,15,17,-62,27,17,12,-4,-24,1,-44,-16,56,1,13,29,-46,-23,-27,-32,2,29,12,-30,33,18,4,-12,-6,20,13,27,58,33,-5,11,-49,-1,3,-32,8,25,50,16,3,-22,8,32,-15,11,26,22,0,16,40,-12,-47,-19,6,-47,32,62,-30,-4,3,35,23,31,57,-25,11,-16,-7,-2,-7,3,41,-16,30,-10,36,40,43,9,17,18,-20,0,29,21,9,6,38,-12,-15,22,-28,-30,-22,-12,-7,30,-23,-4,-43,14,33,19,-1,23,61,4,40,30,-8,-11,-13,-18,-10,-2,29),
	(-2,-34,13,-34,-20,-39,-6,11,-16,16,-38,11,10,14,-13,1,-43,-18,-17,3,20,75,0,0,11,-45,-34,19,8,4,-22,23,-9,-4,-5,-12,35,-15,26,6,13,8,-6,-34,-7,15,-15,23,12,31,-6,-20,4,20,31,-10,5,47,36,14,42,1,-18,-48,-31,18,5,6,17,-2,-30,3,0,18,15,38,-40,23,13,-13,-21,-18,-17,25,-32,24,22,7,-8,0,3,6,-34,-12,31,34,-3,16,-25,40,-22,-6,24,-47,-31,-41,3,29,15,-8,16,-4,-15,12,-18,-11,11,25,-9,43,23,5,-21,-33,0,-23,11,14),
	(-10,-20,-12,-13,-54,-36,-12,-25,10,1,-22,19,-7,6,-65,-8,-17,-7,0,9,1,60,-10,-13,-11,-32,-54,-34,31,2,-34,6,8,-29,-21,-3,2,-4,38,8,9,19,0,-59,-17,28,-26,-12,10,41,10,-21,2,-16,40,23,-23,27,22,12,-6,1,-5,-20,-68,24,-45,-2,26,15,-31,-3,-40,18,25,25,-30,2,6,23,-22,-8,-6,39,-10,12,22,31,12,0,17,24,-59,-8,-9,4,-13,-9,-35,39,-20,3,-5,-10,-14,-22,14,9,39,-13,21,-6,-6,7,24,0,-9,21,-1,26,10,-16,-25,30,1,-18,-12,10),
	(-10,-27,-17,-35,-24,-18,3,1,21,1,-43,-1,9,10,-45,-16,-3,-28,-6,34,8,29,-17,6,7,-20,-48,-12,34,8,-24,5,4,-29,-1,-20,1,-28,20,1,3,13,-32,-56,18,0,-56,-41,17,29,-3,7,29,5,20,39,9,33,37,16,-6,-6,-4,-35,-22,10,-6,-21,50,7,-2,-10,-68,-3,9,41,-6,18,32,4,-26,18,-8,8,0,26,27,35,1,-12,5,22,-31,-18,-20,31,-1,-8,-16,24,-38,-30,10,-23,-19,-19,4,-2,30,-14,21,-1,-19,10,-1,11,18,-4,24,12,25,11,-35,-5,6,-11,7,23),
	(17,-36,-4,-9,-12,-2,3,-15,0,7,-20,19,-13,40,-45,9,0,-10,-10,16,11,49,14,-2,3,-13,-18,-26,8,-19,-20,-7,8,-3,-21,0,19,-9,6,-22,0,23,-67,-70,31,7,-43,-8,6,8,-3,20,12,1,-3,5,-10,7,1,-19,20,19,-16,16,4,0,-6,13,19,-5,13,18,-57,-10,-28,44,5,1,-11,-2,2,-9,2,-20,16,-18,24,-6,4,21,11,37,-22,-18,-28,34,4,0,-3,1,-29,-31,21,35,-2,-1,4,-11,12,-9,24,16,17,15,-6,12,16,23,22,12,36,6,-15,26,-30,0,14,2),
	(-6,-23,-8,8,2,-17,3,19,-20,9,0,46,-35,18,-6,26,-39,14,1,17,-22,10,-12,-6,15,-11,-2,-12,24,15,-27,-22,9,-1,7,-3,-20,17,46,-17,3,24,-90,-40,0,21,-26,2,32,-20,7,16,11,-31,15,19,-7,14,-16,9,4,6,20,10,-21,15,5,-1,27,2,1,19,-41,-30,0,46,4,13,7,0,3,5,-49,-17,26,-18,32,29,-1,4,-16,14,-7,-4,-19,13,50,1,-1,7,-9,-10,20,13,9,-9,21,-24,-13,-9,3,-1,8,29,-7,14,-25,32,31,-4,16,40,-45,-13,12,-11,1,-6),
	(-28,-14,-1,-3,-55,-27,13,8,18,-14,13,21,-36,-9,-3,2,-11,2,0,-3,0,8,6,7,-6,8,19,0,0,8,10,-6,21,-12,9,-6,-27,17,23,-4,29,-10,-52,1,27,1,-37,-14,17,10,23,16,26,-15,-14,-9,23,-1,-5,16,10,-7,-2,-6,-11,-10,1,0,24,4,10,-7,-14,8,-9,24,2,14,11,-12,10,0,-52,-17,6,7,6,6,-24,4,8,34,6,9,-29,12,38,-8,-16,30,-5,-13,21,7,6,3,32,0,16,-11,10,13,10,-4,-7,-9,-4,-2,11,-5,3,3,-28,-37,-12,-23,2,28),
	(-34,-45,35,-11,-19,-34,26,-3,-15,7,-4,37,5,-29,-2,-1,-3,21,-10,4,4,-26,-4,7,7,9,33,-4,16,15,3,7,0,-10,0,1,0,27,0,-6,-5,5,-49,-21,15,11,-15,-13,33,-6,-4,8,25,-5,-2,40,4,7,22,-13,16,-12,35,7,-25,14,11,-1,18,15,5,25,-39,-14,-22,16,3,-2,-8,-9,2,22,-34,19,23,-7,10,-6,-17,11,-22,22,0,-27,-7,17,17,9,1,36,-34,-6,13,36,2,6,33,26,5,-24,34,33,7,3,25,-23,-7,-5,16,-2,14,6,7,-8,-10,-7,14,6),
	(-13,-8,-1,28,-20,-35,10,-2,5,14,20,39,3,-36,6,10,1,17,9,7,26,-27,5,21,10,19,17,-11,11,24,6,-1,39,-16,-9,-14,15,3,-10,7,26,-5,-23,12,26,4,-15,-22,20,-2,10,13,8,-20,-36,-13,36,18,23,-1,37,-1,42,7,-17,14,17,-26,0,-5,-1,28,-16,-5,-12,-24,2,-5,-23,12,-21,7,-42,17,26,-19,39,4,4,0,-43,11,-12,-22,-5,1,20,13,-12,-8,-33,14,8,10,41,14,-1,28,-28,1,14,29,32,9,-2,16,19,3,24,-5,9,10,-10,-9,-23,25,28,10),
	(11,0,7,29,-21,-35,16,19,-9,27,21,71,-30,-46,3,24,-23,15,30,17,6,4,-28,41,38,-19,47,-11,11,24,8,-33,27,-8,8,6,-3,24,-5,15,-1,-13,-6,-15,23,13,-13,-12,34,23,0,20,7,-1,0,-8,18,2,6,-8,8,-12,23,-21,-4,20,-9,-17,9,24,-2,30,0,-6,-31,-12,-13,17,-21,1,3,16,-38,-1,16,0,31,11,13,-21,-15,28,-4,-19,-4,18,14,17,-25,-29,-38,1,15,5,29,13,4,4,-20,-4,-9,19,32,18,31,-18,3,-11,-3,22,28,27,2,-15,-12,4,11,9),
	(14,36,-2,13,-4,-41,4,27,-4,17,33,56,-10,-2,-16,39,-26,14,36,16,-23,0,-15,12,31,-6,26,13,13,22,4,-15,32,-1,26,13,-5,8,-15,28,-4,15,-3,-14,33,-1,4,-4,15,18,16,19,-6,-30,-4,7,-4,0,6,0,3,26,8,0,1,-8,-41,-19,28,11,13,20,-24,18,-42,-6,11,6,-25,0,14,3,-31,-9,35,-7,49,14,20,1,5,18,3,-25,-10,7,14,27,-15,-43,-10,2,-7,2,-1,21,0,31,-47,-8,0,3,12,31,23,-19,12,27,6,16,29,-18,-4,16,-27,21,9,-7),
	(-3,38,17,21,-11,-18,-1,16,-14,16,4,28,10,-33,-7,24,-41,0,19,11,-7,-4,30,1,15,14,19,5,-2,4,11,-15,5,9,0,-10,-10,0,26,14,15,-2,-2,6,16,-39,8,0,24,-3,10,10,-5,8,-30,-20,25,5,-5,3,-12,-6,-11,-8,9,4,-47,-10,10,12,-3,19,0,-15,-16,12,0,-7,-18,-7,22,6,-43,-19,16,-38,17,-13,18,4,10,3,11,-26,18,13,-4,1,-51,-42,-21,2,-23,1,21,28,-8,20,-29,12,23,15,32,13,12,-6,31,-11,-9,8,29,-20,4,5,-12,13,35,-7),
	(13,37,-1,19,2,7,-17,23,2,1,6,42,0,-27,39,17,-23,-1,21,0,-10,21,0,-6,-3,26,21,14,7,-19,10,-3,49,-22,1,8,-8,-21,23,22,13,-14,2,-15,28,-43,-4,-12,17,20,-16,9,-10,-11,-35,17,34,14,-6,17,-17,4,-27,-6,12,33,-29,-14,1,-5,12,-8,-9,6,16,-3,-2,8,13,18,3,29,-57,-30,21,-2,31,-17,53,-7,-10,1,4,-37,-5,-24,-6,46,-28,-56,-27,30,9,30,-23,5,0,53,0,29,7,0,11,16,23,-11,46,-5,-8,11,15,-11,-28,27,-32,17,33,-11),
	(-8,36,6,10,27,-14,-20,42,0,36,32,29,12,-25,12,24,-18,0,-8,4,12,41,19,-67,-14,9,-5,-1,7,7,21,-10,44,-4,-1,-7,0,-27,0,31,14,-46,13,4,11,-7,-5,-30,7,11,-37,18,-31,19,-13,0,-1,5,-28,-10,-16,21,-36,1,0,-9,-31,-22,20,11,3,13,17,4,2,-3,17,5,-20,-15,14,37,-75,-25,12,0,9,-4,0,3,20,20,6,-2,-1,-29,-4,29,-29,-66,-41,7,-21,-9,-36,15,-14,15,-18,21,-18,9,-3,-22,-4,8,4,15,-10,17,9,-13,-6,6,-18,15,18,18),
	(5,32,22,43,35,11,-26,5,-12,30,35,16,9,-12,13,27,-43,5,-20,13,-19,46,-11,-63,-8,53,-12,-6,-8,-15,57,-28,12,16,13,10,7,5,23,7,2,-49,-9,38,39,10,-24,6,-4,-38,-22,33,0,2,-26,0,-27,-6,-55,-4,-23,1,-33,20,2,-23,-42,7,-20,3,35,-6,15,-21,23,13,27,29,-22,-35,35,48,-46,-56,16,-21,-10,10,18,1,-29,-2,-22,-42,-7,-22,0,28,-24,-40,-13,0,-22,13,-6,20,18,0,10,-13,14,28,-3,-1,-49,2,-7,0,8,-17,36,3,23,38,-8,14,45,1),
	(-26,8,-1,37,19,-16,-16,12,7,-4,42,12,6,0,7,15,-19,10,29,-24,2,49,-29,-25,11,26,4,-7,-32,-16,31,-21,-4,-34,22,18,15,19,13,-21,-1,-37,-8,31,16,-10,-2,-20,-17,-16,-48,27,9,12,-6,29,-15,-21,-18,-3,-34,-5,-48,-8,-18,6,-42,-30,-15,5,6,-14,-1,-21,23,-17,32,7,-14,-22,3,10,-66,-44,-2,3,19,-34,1,-27,8,-6,24,-28,17,-15,5,26,17,-33,2,37,-10,36,12,17,19,-3,-27,-4,9,8,9,19,-33,-28,-21,-33,-21,-5,19,-6,12,38,-34,30,34,17),
	(-21,36,18,11,12,-5,18,44,14,4,18,5,6,17,16,20,-22,-13,-6,-27,-20,24,-28,-9,17,41,-5,11,-27,-4,33,3,15,-20,3,12,-15,-7,4,-26,-16,-11,-28,4,36,12,2,-25,-23,-10,-23,2,-25,12,-24,22,-24,-1,8,-9,-19,5,-43,-21,-41,26,-28,-21,20,-23,8,-10,-9,-25,36,-14,22,28,17,-17,13,28,-28,-35,-19,23,-17,-23,-19,-31,2,-6,18,-44,24,-28,4,48,9,-3,-3,-6,-43,17,-19,-26,35,-3,1,-13,38,24,0,-17,-19,-24,10,-20,0,-7,-5,-15,13,10,-15,19,7,43),
	(-8,10,19,12,37,10,-21,31,26,1,3,-23,24,23,0,-1,1,27,-10,-22,-33,1,-23,-5,-30,38,3,27,-11,10,12,-10,0,-16,-16,23,0,28,-19,0,16,-9,20,30,29,4,5,-18,1,-37,-27,24,-8,25,17,20,-33,-7,-25,-15,-30,20,-2,7,0,-8,-41,-17,18,27,36,5,-29,-12,-13,10,8,2,13,-16,-1,27,-16,0,1,0,-7,1,-20,-6,-10,-10,-14,-14,2,-32,-41,34,20,19,-9,-8,-24,11,10,5,4,-14,-8,-32,25,21,2,-12,18,-25,-3,-31,-14,3,4,-41,-15,27,0,0,0,8),
	(4,10,24,11,-9,9,-12,23,-19,-22,11,-14,-11,27,-21,-5,-7,-15,-17,-19,-36,-26,-21,7,10,47,26,20,-8,0,23,-5,36,-12,-16,4,-4,-1,1,-17,-35,-6,-20,-2,59,2,-36,-44,-20,-19,-23,8,-30,28,4,13,-13,-34,-13,-7,-35,-4,-20,0,21,-5,-17,-21,0,-11,26,-28,-45,16,1,-11,34,12,13,0,24,37,-48,-16,-15,8,-4,27,-2,-12,-11,2,-2,-1,-3,-15,-37,22,33,23,-9,-5,-5,21,-17,-5,2,-6,-3,0,24,20,-10,-6,4,-12,-3,-45,12,-30,-12,11,-9,20,-31,-9,1,3),
	(31,32,36,26,-19,0,-9,37,-4,-46,29,-13,6,37,-20,10,-17,-8,-9,-17,8,-22,-5,23,23,7,-14,15,-15,-11,27,-25,30,-28,-6,-2,-15,-2,16,-28,-6,-15,3,15,36,-1,-53,-9,-23,2,-26,5,-40,45,-5,-9,22,-19,8,16,-23,17,-10,3,34,10,-31,0,14,-11,36,-46,-35,-14,-12,3,40,30,0,-48,38,50,-7,-27,19,-6,22,-8,0,-29,10,17,12,-27,11,27,-31,58,34,-16,18,-22,-30,-15,-10,-27,18,-49,1,-31,9,59,13,-53,-11,0,4,-29,39,-17,-29,6,18,0,-55,13,-32,17),
	(20,-13,-9,6,0,13,25,-8,-9,-3,14,-22,21,20,-35,34,-14,26,-15,7,2,-3,32,-2,6,0,-1,63,9,-7,27,-19,24,-15,-4,-42,24,15,-22,6,7,-15,21,3,-21,-9,-30,-20,-30,-11,7,3,-1,20,10,-20,-8,7,-6,17,-10,13,-6,-24,26,-18,-36,5,19,-21,26,-17,-23,1,9,36,23,26,5,-34,-7,7,-4,-52,32,-24,9,13,-19,-29,-15,15,2,0,-20,13,-10,51,3,0,23,-44,-12,-19,-26,-21,-8,-31,-40,-14,0,57,-30,-32,-52,-13,-13,15,-8,1,28,19,11,52,-32,8,31,-20),
	(-4,-23,-9,14,-10,7,0,15,6,9,15,-20,31,0,0,27,24,-5,-18,7,-28,-7,-2,-9,-7,12,-13,0,-12,33,7,-14,22,-35,5,17,0,-6,6,2,-38,-12,19,14,18,-11,-6,-5,-40,-7,-17,9,-23,-10,34,28,-4,12,-1,4,-32,20,22,20,-23,-4,-25,5,15,-16,-2,7,-20,8,-26,4,6,3,0,-2,-9,4,15,-3,-1,9,5,23,-2,9,10,-6,-21,20,0,-7,-9,1,20,-3,23,-4,-13,-15,-5,10,-10,-32,-22,-9,-27,6,10,-9,1,-24,-12,-31,-16,3,2,5,31,8,0,-14,27,-16),
	(1,3,-21,-2,16,-2,-1,2,16,-9,19,-42,1,-13,10,15,10,19,-13,23,8,15,19,-16,-10,-8,15,-3,15,19,19,-16,-15,10,-4,14,1,15,2,-25,-4,-17,-7,19,-3,26,18,4,-31,-1,-15,3,5,-5,-5,22,-5,-13,-1,7,3,-3,15,-24,0,7,-24,-9,-12,-3,0,24,21,0,-22,18,6,-9,-9,12,-2,-26,27,14,14,13,19,18,6,33,7,-13,-19,4,-6,-12,-15,0,11,15,-5,-1,-21,23,20,8,-11,13,0,1,-11,16,-1,-2,-6,-1,-8,31,8,17,-6,23,28,13,19,-13,-9,5),
	(7,-4,17,-11,-19,8,20,12,-1,8,0,9,-13,-1,9,8,-18,9,10,13,-8,-9,16,9,-3,3,12,6,12,-5,14,-19,-15,11,6,-6,-15,-4,8,-8,-8,18,18,19,-8,10,-7,-10,17,-9,-3,-10,-17,15,1,0,19,-6,-1,17,-16,16,-4,12,0,0,-18,-13,-7,-9,-19,-3,-3,13,-7,-18,9,-13,16,3,-13,9,6,15,-20,-15,-6,-17,12,-13,-5,11,2,14,-10,-20,-9,19,-15,11,-9,7,-1,-18,-20,-15,2,12,-19,-3,-10,-4,-8,-12,-19,-20,-18,7,12,-16,-2,-7,15,10,6,15,15,-4),
	(-9,-10,3,-16,2,-19,-16,18,6,-4,20,5,-20,-12,-19,-20,-10,11,-15,-15,-1,0,-7,15,15,6,-18,16,-15,-8,18,-3,-4,12,-8,-20,-12,-6,17,-6,8,-4,15,0,8,-3,11,12,17,5,3,-6,15,1,5,2,-19,14,20,-3,-3,14,-16,-15,5,-6,-15,15,0,-10,-10,20,11,10,8,-4,13,4,-14,15,-16,3,2,2,-6,8,-8,1,0,2,-1,18,-3,9,-17,-6,-18,-8,-5,0,17,-20,1,-16,-11,15,2,20,-5,-16,20,-18,-10,18,-9,12,9,-19,9,-2,-8,3,-3,-7,6,-6,-20,-18),
	(-7,15,-3,2,-17,-2,19,9,20,-13,-2,2,-17,-17,10,-9,-13,4,-10,18,-13,19,-2,-8,9,6,20,-1,15,19,2,-6,0,16,-8,20,2,17,-14,7,4,-2,20,-18,0,-18,17,13,19,-12,12,-14,-2,-8,-1,-15,-19,16,17,12,-10,0,-15,1,-11,10,-19,4,-14,-8,14,4,-18,-4,-7,18,0,-13,-14,-3,-17,17,-1,-14,3,-11,8,20,6,2,-3,-1,11,-1,11,2,-17,-1,-6,-16,-18,-16,15,-9,5,1,9,-2,2,3,0,17,-9,3,-11,-13,12,6,-17,-7,12,17,3,6,20,-6,8,2),
	(20,3,2,19,-25,17,-15,6,-8,8,-22,3,4,23,-25,-14,12,-39,-7,10,-18,-19,-18,16,-5,12,-23,40,-21,-16,-1,25,9,3,-3,4,-30,11,14,-21,-23,0,3,4,29,2,-6,-42,-37,11,-11,19,0,19,-6,-15,11,10,6,12,36,22,-19,-1,6,-9,11,8,-4,-12,5,7,14,1,0,19,-16,9,-32,-6,13,-1,11,-30,30,-15,-31,0,7,19,-13,34,3,-2,-22,13,17,17,5,-11,7,9,0,15,-28,-19,3,-3,-6,-6,10,23,3,-26,7,6,17,0,20,28,-16,-10,9,-9,-1,20,-42,11),
	(35,-17,37,-21,4,-12,24,0,-18,-24,-41,16,14,9,-4,5,19,-4,24,9,19,29,33,3,5,-12,2,-24,2,26,9,-12,-27,0,16,-20,2,-27,22,-4,35,9,12,-15,-22,0,28,14,7,4,0,-15,9,-2,16,-8,31,-2,17,2,-11,26,25,-19,0,14,0,-6,9,26,-24,-7,-1,-24,-10,-11,19,-36,17,-12,-1,-12,-17,8,-3,21,14,-12,-32,21,-9,-7,12,-5,2,-25,-4,12,15,10,-24,33,-6,-28,24,-17,2,2,5,15,1,9,1,8,-7,-24,-26,8,-19,-15,16,-3,-3,-38,31,10,40,-16),
	(-34,-19,13,-47,-35,-17,5,3,-18,20,-18,-8,9,51,-16,-28,13,-18,3,41,-6,37,47,-20,26,-15,-19,-23,12,10,-12,37,16,18,16,-23,25,-38,0,32,18,3,11,-39,5,-6,-38,-11,18,29,-35,-32,-1,11,49,11,24,31,-2,-5,11,20,-2,-48,12,2,-30,-20,30,9,-20,-22,26,13,-11,14,-32,16,24,13,-30,-9,-2,41,-49,23,1,23,9,20,5,-13,1,35,4,-3,-3,55,14,16,-14,0,6,-44,3,-52,11,25,34,21,6,-2,-42,0,-22,-2,-19,36,-6,-4,21,-18,23,-20,28,-12,-4,14),
	(-10,-21,23,-30,-35,-5,11,-25,18,-12,-24,-14,-20,22,-45,-62,-27,-51,-38,8,-30,44,8,-42,6,-29,-65,-15,19,2,-20,26,37,-10,-13,-39,11,-24,47,23,-24,-7,44,-24,-12,21,-41,-15,-11,55,-31,-19,-11,23,41,28,29,14,18,18,23,26,1,-49,-17,-18,-24,-12,50,1,4,-19,46,33,37,49,-4,23,11,-13,-17,17,28,12,-34,37,-20,25,8,22,2,24,8,24,23,17,2,32,-14,34,2,5,29,-50,-57,-47,18,0,58,17,-8,-15,-34,10,28,-2,-1,4,5,13,10,-16,-18,-41,22,-28,-15,68),
	(-7,-18,11,1,-48,-9,-2,-36,47,15,-1,12,1,5,-27,-41,-25,-19,-6,40,-36,17,-33,-7,-11,-13,-61,9,34,-1,-5,43,37,0,-15,-30,-4,18,-20,-6,-30,1,-10,-68,24,35,17,-29,20,46,-44,8,0,0,40,-8,-6,25,-5,16,43,14,-26,-25,-33,-27,-62,-1,40,-11,11,25,14,-4,55,7,3,0,17,-6,-20,1,-8,-46,12,-21,4,8,19,19,-21,25,-4,-16,-3,17,23,32,-9,33,11,-2,37,-5,-11,-22,10,3,23,-26,-12,-12,-7,47,16,26,7,23,-23,17,8,-9,-25,4,9,13,-22,36),
	(10,-8,0,-11,-40,-21,-16,-31,44,14,6,31,9,2,-40,-26,-56,-24,31,25,-12,-3,-19,-25,5,-15,-67,21,19,4,-9,22,25,9,-17,0,-20,-14,-12,8,16,5,-45,-51,-4,-3,-36,-28,4,19,-33,-2,6,18,24,13,-5,47,1,9,33,0,-7,-19,-23,-6,-29,2,55,4,-6,15,14,27,38,5,-15,-1,0,-12,-23,0,-9,-19,15,-9,24,19,8,35,-36,7,-35,-6,5,27,0,44,-24,5,-15,-33,30,-28,-3,-26,8,33,20,-46,25,-26,17,9,16,-5,22,24,-19,37,24,-8,13,-6,-13,-21,0,5),
	(1,21,-19,19,-7,-18,-10,-19,48,3,-4,30,-24,13,-11,-20,-17,-27,20,28,-9,-23,8,-27,-26,-15,-51,34,12,9,-28,44,30,0,-47,8,-4,-12,-8,25,38,-2,-53,-39,-6,7,-43,-31,13,41,-28,-9,14,22,28,-5,24,45,2,-15,25,43,-3,-12,4,-35,-15,-18,81,-24,17,22,-8,18,62,10,-30,18,-7,-25,-10,-11,11,-12,-8,-7,13,28,-6,16,-32,38,-48,-10,-9,2,-4,23,-36,23,-21,-15,9,-17,-37,-33,29,1,17,-36,27,-37,-20,7,41,20,23,38,7,49,37,-45,9,11,-43,-10,16,21),
	(-6,15,12,-3,-47,-23,-11,-32,-5,6,-20,25,-44,8,-11,-4,-30,7,11,1,-10,-47,-14,-13,4,-11,-25,4,2,-11,-20,23,16,-4,-17,-13,-1,7,18,26,40,19,-93,-45,23,33,-10,-20,31,43,-4,-31,28,0,0,24,51,33,22,-6,48,16,4,6,-1,-18,-12,-15,47,-15,-2,27,-27,8,27,7,-29,21,5,-25,-30,8,-45,-15,-8,-14,-17,15,16,24,0,23,-30,-31,-8,7,9,38,19,48,-6,-35,39,-6,0,-33,23,-6,26,-29,33,-10,16,29,13,0,7,27,-7,40,30,-36,-13,-4,-17,5,28,38),
	(7,30,6,-9,-90,-23,40,-40,23,-8,-37,39,-50,-15,-18,-4,-29,-25,20,-3,0,-40,-51,19,-2,21,-31,15,-9,-4,-31,-1,49,0,5,5,-4,5,-3,12,-6,9,-86,-45,7,10,-5,-21,35,42,-29,-12,6,35,20,7,42,47,30,-19,33,27,18,2,0,28,-20,-5,46,0,6,12,-29,4,1,6,13,19,9,-8,-40,12,-50,0,-25,-11,3,-21,-4,20,-32,2,-23,-63,-7,4,-20,78,-20,47,-7,-22,20,-22,-22,-33,8,52,-6,-14,28,-32,37,46,37,0,9,0,-12,36,8,8,-35,-54,7,-10,-1,12),
	(6,4,46,-2,-67,-21,6,-34,-10,-17,-47,24,-16,-17,14,-20,-35,3,26,-13,-15,-19,-57,-11,26,-14,-5,10,-9,-15,0,17,51,-4,-8,-22,23,-4,3,34,14,-1,-90,-41,-8,32,-27,3,46,45,-8,-34,8,-2,-7,22,37,12,35,-2,30,35,15,4,-34,13,-30,-26,25,3,15,18,-14,13,25,-21,-17,18,1,-3,-16,20,10,-12,-35,-11,0,-20,-21,10,0,25,-23,-28,12,4,-18,58,-36,52,-10,-16,28,-11,21,-21,21,36,-24,0,23,-33,-10,13,45,-2,20,7,5,33,11,-7,-7,-28,0,1,33,43),
	(11,-5,17,24,-58,-26,17,6,20,10,15,30,-18,-22,-6,-1,-20,-23,21,-2,14,-19,-78,-19,10,23,4,31,15,-6,21,26,34,-10,-29,-3,7,0,-7,38,24,-2,-56,-26,-12,26,-27,-20,27,22,-19,-18,14,4,22,-12,40,25,-17,8,40,26,1,-5,-16,-20,-11,-23,53,2,9,14,-9,27,13,0,-15,4,-22,-20,-20,15,-22,3,26,9,34,18,5,9,-30,-12,-33,-45,1,30,-42,34,-68,8,8,-36,5,-11,-1,-33,4,30,-12,-49,-9,-23,-12,18,3,13,4,35,-8,56,43,1,0,5,1,2,11,6),
	(4,28,17,3,-19,1,24,19,15,10,-18,58,-15,-6,-11,-30,-41,-30,-1,4,-12,5,-67,-36,-3,18,0,30,8,-31,42,45,15,11,-10,-3,20,6,9,14,1,-28,-33,-39,9,13,-46,-6,39,17,-1,9,12,13,24,5,45,31,8,-16,39,10,19,-8,-9,-12,-24,-22,48,5,32,6,-14,19,5,2,-10,23,5,-24,-35,9,18,7,17,-15,16,47,10,-8,-10,-21,-40,-17,13,3,-23,51,-104,-21,-17,14,7,9,9,3,8,-8,-7,-15,-3,-32,-1,38,36,7,32,17,-26,23,36,-5,-12,-25,-11,18,12,37),
	(27,16,0,20,-33,4,0,40,27,-1,26,26,31,-20,2,-24,-50,13,3,2,24,9,-34,16,26,16,17,-1,-5,-39,48,40,-7,5,10,17,2,17,-17,2,-8,-13,-9,-12,-8,9,-69,-6,10,24,17,-28,24,5,-1,38,11,-14,-4,10,24,16,-4,5,3,6,-43,-36,14,-11,-2,8,-7,7,0,-6,15,12,24,-14,-39,30,4,0,0,-5,40,35,-2,-17,-7,-6,-11,-21,34,23,13,35,-113,-39,-8,9,13,9,6,-5,25,42,-15,25,41,-18,11,14,39,15,28,-22,8,6,22,-12,4,30,-10,8,-6,6),
	(-2,-18,20,7,-23,-6,-19,52,20,-7,9,33,24,-44,23,20,-30,21,4,14,27,2,-10,-33,12,5,2,23,-1,-47,43,9,10,-1,-7,-11,11,-10,8,-7,3,-8,3,-11,-5,-34,-47,47,3,1,22,-9,11,6,-9,7,20,0,-4,-13,30,4,6,-25,-19,17,-24,-16,37,-9,10,12,16,-33,-15,7,19,-17,3,11,-16,24,-4,0,4,-11,38,3,7,-15,-27,16,-10,-29,7,17,23,60,-74,-21,-7,23,18,0,-12,17,16,30,-44,-7,13,-22,14,15,45,-30,4,5,1,33,65,-27,-4,12,-5,18,56,6),
	(-3,9,-14,28,-49,-8,-8,51,20,-8,12,34,18,3,15,20,-17,6,1,-7,15,20,-30,-57,37,23,15,15,-46,-60,29,27,34,-14,-21,-18,9,-33,-12,-4,27,-57,-13,-20,-6,-53,-38,16,21,4,29,0,4,7,-12,20,4,-7,-11,2,40,5,-9,-26,-16,3,-36,0,37,15,0,1,52,-28,14,17,14,4,11,-18,-18,3,11,-36,-9,-5,20,10,-5,-30,-47,-1,-7,-59,-8,19,7,69,-57,-28,-32,4,16,-11,-13,13,13,29,10,12,31,-36,-2,4,25,-5,30,-8,8,26,58,-43,4,16,-20,37,18,-3),
	(6,-11,31,7,-19,-12,-16,18,-1,-5,-10,0,21,9,-5,26,0,26,32,19,17,51,-12,-40,24,10,-4,-1,-20,-19,37,3,54,18,4,25,10,-16,25,-11,33,-29,13,-1,28,-37,-30,13,-3,17,-7,14,-3,27,-12,22,37,-35,-30,-22,-14,39,-22,-15,38,23,3,0,37,0,10,5,49,1,19,11,31,10,5,-41,-13,19,-26,-14,-26,-11,38,-29,22,-28,-10,8,27,-50,16,15,-9,63,-15,-29,-32,37,-11,19,-14,13,1,32,-15,1,-1,-41,9,5,-8,-13,15,3,-3,35,52,-27,-2,23,-32,33,22,8),
	(6,14,17,3,23,-24,-7,-5,9,-13,-25,-16,23,-4,24,1,-6,-12,17,4,22,51,-27,-40,13,24,-2,8,1,-5,28,-8,14,15,-8,20,-2,10,26,-19,10,0,-27,6,14,-20,-31,-1,-4,2,-7,7,9,36,1,3,26,-14,-19,8,-36,-16,-54,-10,-1,16,-15,17,44,-28,25,5,-1,-15,13,24,22,14,-16,-47,-11,13,-34,-25,-16,-6,29,-15,-7,-3,-39,-12,4,-50,-14,-5,-2,52,5,-7,-3,8,-38,-12,18,1,-6,13,-6,15,-1,-29,12,-1,-29,-44,26,0,3,20,41,-45,9,32,-26,1,46,30),
	(11,4,15,4,-18,-51,20,24,0,14,4,15,-11,8,3,-17,-44,-15,15,-4,13,68,-23,-1,41,30,-40,6,-9,-14,46,19,51,-5,-12,11,17,-10,0,-6,23,-1,3,-23,-9,-10,-25,-28,10,0,-29,-23,19,53,10,-17,21,13,-2,-16,-5,-40,-67,-27,-20,25,-5,4,34,3,12,-2,42,25,39,2,6,25,-42,-74,-1,16,-48,-39,2,-35,22,-4,-12,0,-31,2,5,-36,-12,-6,-1,70,51,-8,-10,10,11,-16,7,3,-10,20,3,-16,19,-10,3,37,-16,24,26,23,9,52,36,-16,-1,11,-59,6,-16,28),
	(33,50,30,32,-7,-19,8,6,17,11,-24,12,2,28,-19,-24,-63,-32,6,-47,6,35,-43,17,19,16,-14,34,-7,-10,38,13,55,0,2,4,6,-3,-25,-14,4,0,-17,-15,-3,-20,-10,-27,9,-7,-45,-27,-24,36,-6,-19,-16,-1,-19,18,4,-8,-37,-18,-7,9,-37,-18,15,-3,33,-9,35,3,26,30,0,41,-10,-44,-6,51,-46,-66,6,-13,39,-4,-18,-3,-15,0,-14,-22,-1,-18,-21,71,24,-6,21,20,10,12,-14,-2,14,-10,-18,-44,8,32,11,-7,-23,42,19,0,-13,10,19,-22,-5,-16,-44,22,-8,15),
	(21,25,35,21,-15,-23,-3,16,-42,29,-38,5,-6,50,0,-8,-50,-12,-9,-23,10,6,-22,-13,44,0,-23,23,-44,14,10,20,13,-11,4,13,35,-9,17,-11,0,8,-41,1,-3,-17,-51,-22,10,-39,-23,-27,8,25,-15,4,-9,-13,-17,-4,12,-20,-31,-29,-17,33,-27,-18,33,12,-4,-17,44,-3,18,-10,34,4,-20,-35,-16,10,-50,-51,-31,-8,28,-14,-27,-21,26,-4,34,-31,3,-25,-12,14,39,5,9,-20,-29,-22,-23,-14,35,-8,13,-6,35,3,-5,12,-64,-8,16,-5,-3,-13,26,-14,-1,21,-19,15,-9,44),
	(34,16,69,-19,-23,3,-8,4,-48,25,-6,34,-24,44,-6,-19,-25,-15,-20,-28,13,21,-62,-1,35,-17,-6,-7,8,-19,8,3,-6,31,9,-23,50,2,24,13,0,38,-49,-51,31,9,-18,10,18,-22,12,1,17,22,-29,-34,15,-18,-25,18,15,-17,-11,-18,-6,45,-43,-17,34,19,2,-14,14,-23,12,13,31,15,-15,-39,22,6,-46,-46,5,5,21,37,-34,9,29,2,29,-20,-19,-9,-17,-8,25,9,0,8,-33,-28,-17,-24,-25,-22,8,-31,5,35,9,12,-52,-18,10,-23,-6,8,42,23,-22,-1,-14,37,-8,19),
	(51,19,39,17,23,0,-18,14,-49,-24,-28,31,-43,34,-18,9,12,-17,-6,-25,22,-44,2,34,10,-34,18,-2,2,-13,31,-12,-6,4,17,-22,9,22,37,26,37,13,-37,-42,25,-5,-33,0,12,-19,-13,13,9,3,-18,-10,15,-14,-11,-2,-20,-7,-35,-34,14,33,-29,7,28,-6,-30,-11,-6,-42,-29,13,59,-2,-26,-17,57,38,-10,-8,-8,1,29,40,0,-26,25,-3,13,-2,-26,5,-39,17,-12,10,26,-9,-20,2,-25,-45,2,-12,0,-4,-33,41,9,-8,-48,20,-10,-33,45,-1,-10,5,-7,-39,-12,7,-24,2),
	(29,4,28,-3,15,-27,-2,0,-21,15,-3,29,-24,34,-34,7,-16,39,-4,15,21,-18,24,-18,20,-12,30,12,-5,12,10,-3,24,17,-15,-41,17,23,33,25,24,9,-7,-47,8,-4,-1,-7,0,1,4,1,30,19,-10,-27,0,-13,0,15,-15,-17,-32,-36,4,22,-14,1,10,3,0,13,-17,-36,21,39,10,-3,-37,-27,1,-4,-4,-2,6,-19,26,24,9,6,17,12,8,-18,-10,-12,19,19,1,10,14,-26,-24,-7,-14,-45,-5,-16,-17,-4,-20,19,-2,-3,-56,0,-12,-3,15,17,29,27,-20,-5,-20,22,-2,-18),
	(-18,-18,-6,14,0,13,19,3,-1,-9,10,-36,-1,-14,20,5,11,-9,1,1,-20,-15,4,9,-12,14,-8,28,-4,-6,-5,6,26,-2,12,2,1,-18,-2,-11,-18,-1,7,9,5,18,-13,6,-35,-6,-1,-8,-19,0,-4,33,8,-1,11,-9,4,5,9,0,12,7,10,-19,-1,4,12,8,-16,12,14,29,-2,31,16,-16,-3,17,7,7,7,-1,17,22,-14,20,-11,-13,-1,-13,0,0,-9,12,16,-15,10,7,1,3,15,-8,6,4,3,1,-16,24,-6,-4,-12,-18,13,-2,12,22,-10,8,10,-17,-4,-3,-16,-8),
	(-21,-33,-26,28,0,2,9,0,26,-3,10,0,-10,-14,-10,-6,2,18,5,7,-24,8,-7,11,13,22,22,-6,2,-17,1,-16,13,-2,2,5,23,11,-7,-9,20,-14,28,18,-25,-20,24,8,-1,-11,-14,-7,14,3,23,0,12,-12,-2,-9,-9,15,-8,-24,-7,-10,5,17,12,-20,8,27,15,-3,-26,16,5,13,-23,0,-15,1,26,-1,-12,-2,-11,10,8,11,12,1,13,8,-8,-7,0,-17,13,-13,14,-17,-17,20,23,12,-12,2,-7,-3,-12,-9,-1,0,10,11,0,-18,-15,19,24,9,24,11,17,-10,2,-8),
	(-11,17,13,10,8,1,-13,-18,3,-20,-16,2,3,10,-14,5,-2,-7,-15,-1,7,-7,13,-12,-16,-11,0,3,-7,-17,12,-9,19,17,-19,-14,0,-16,11,-20,5,-15,7,8,18,11,4,-16,20,0,-15,4,14,4,2,-16,-17,-19,-12,4,16,10,16,16,-9,16,-7,-13,8,-8,11,7,-19,-18,-1,14,-16,-2,-8,2,17,18,-18,4,-8,1,0,0,-12,6,-6,-11,11,11,3,0,-2,17,-5,0,8,-19,11,0,19,0,-11,15,13,3,-14,-11,-13,0,-20,0,15,-18,12,-3,-13,-14,-8,10,13,-17,16,-1),
	(-8,-9,7,3,17,-5,-4,-6,19,19,-11,0,17,-9,-11,-1,8,-2,17,-6,17,13,-3,14,10,15,-7,6,-19,-17,-1,3,-6,18,-12,-7,1,4,-7,19,-18,10,-7,-11,-9,-4,-13,6,4,-15,-13,-7,8,12,15,8,-6,8,-8,-17,4,9,6,-12,-2,-5,-12,15,-3,-6,7,8,20,-19,-15,12,10,2,-4,20,-17,-4,18,-10,18,-5,-9,18,-19,-19,20,4,1,1,11,-8,1,8,-17,-8,-17,-10,-15,15,7,10,17,-16,17,10,-13,-15,1,-1,-19,5,16,-7,-13,16,18,3,11,7,14,-11,-1,12),
	(-5,16,-11,-14,5,1,3,15,-13,19,-18,8,-2,-4,8,-18,-11,18,-6,-7,-13,11,-12,17,-15,6,11,-5,-17,7,-19,8,-17,-12,15,10,-11,16,18,18,0,10,0,-12,1,10,-7,0,-13,8,10,-17,-19,-1,4,6,-17,12,-9,-1,18,15,-15,-12,11,-6,11,19,-10,-9,-15,4,-3,-13,12,-8,-15,8,10,13,-14,13,18,8,-15,-12,-12,0,2,18,-7,5,-1,-7,6,-5,10,-10,14,10,-2,-7,-13,17,14,18,4,-18,17,-5,1,-15,6,-9,4,-18,8,-18,-9,20,-3,-5,6,8,-19,7,-1,-3),
	(12,-2,-11,18,-4,-9,10,-5,-17,5,-7,2,-14,-15,0,-2,5,13,11,3,-1,-4,-4,8,10,12,11,8,3,20,-8,-16,0,-1,6,-17,13,17,-15,6,-11,7,-1,13,-12,-11,-8,8,-12,-3,13,18,19,-12,0,-14,9,3,19,-6,4,-11,18,-20,17,18,-15,-14,-6,2,-2,-15,15,2,4,11,5,-7,-10,-2,-18,-10,-3,9,-1,14,-2,20,6,11,-11,-1,19,15,-7,-17,-11,17,-2,-15,-17,18,7,2,20,7,11,-14,-16,2,-4,-7,-10,-14,3,16,-19,0,15,-6,-2,-20,11,-1,-13,-17,-10,13),
	(-7,-15,3,-5,-5,-16,24,-3,-6,-17,-9,-20,14,-10,6,14,-3,-8,14,9,8,7,-17,8,-8,-18,0,24,-22,-2,6,23,-9,-6,6,16,-2,2,-9,6,0,-1,7,17,15,2,-25,16,15,9,-11,-9,-17,0,12,-11,6,-2,-14,-14,1,11,-23,-2,21,-2,16,-7,9,-8,9,-21,27,3,10,22,-8,-2,-17,0,19,14,-5,2,-12,2,-4,14,3,7,6,25,0,8,6,-1,-11,19,2,-26,4,1,-5,-20,-4,-19,10,3,12,0,-10,1,-9,-6,-7,9,-14,7,7,3,-5,18,8,18,-7,22,3,-14),
	(27,19,20,-10,11,47,19,10,-12,-15,-4,-3,-44,-8,-4,-31,-1,-41,-30,0,-43,6,14,24,-11,45,-23,-8,5,0,31,0,-3,1,-5,-3,-23,-17,10,1,3,-29,14,30,32,3,-25,4,-35,-4,-23,27,-52,-17,-31,40,39,-35,-22,-4,12,-4,-19,27,38,7,7,37,29,-16,39,-22,6,-27,-5,16,35,17,-17,-21,32,48,31,-22,15,9,-17,-16,32,-17,-14,38,22,22,4,25,-2,9,-5,-25,16,2,26,-10,-32,-3,16,-21,34,-1,-1,22,6,-25,10,0,11,-20,21,-41,0,14,29,-41,-18,-14,-28,29),
	(39,11,22,-7,-6,2,-22,-4,-18,4,-8,16,-31,11,-10,-42,-10,-31,-17,-11,-10,9,20,1,-15,10,-34,0,-31,-28,19,4,45,4,-25,-21,-35,4,23,-18,-40,3,16,3,42,1,-34,-8,-18,-17,-50,-6,-41,28,11,35,37,-6,1,1,-4,-16,-68,-17,-21,-26,-13,15,-39,-46,41,-55,-1,-6,9,8,21,25,-9,-36,1,56,14,-54,0,4,3,-1,-3,0,-18,43,15,35,-8,24,8,37,-17,0,34,7,33,-22,-66,0,25,-7,37,-5,9,21,-10,-34,-13,21,7,-45,49,-40,-16,21,-11,-20,-3,17,-48,54),
	(45,13,19,-16,-15,-10,-4,-3,-4,3,-11,0,-11,31,-6,-48,-34,-65,-16,-21,1,26,13,-10,-2,0,-34,-24,-14,-11,7,40,14,15,-27,-39,-12,-22,12,0,-15,7,13,7,25,-17,-59,-15,-33,26,-79,-1,-43,20,2,13,36,-6,-10,16,18,11,-36,-6,14,-7,-17,17,-38,-27,16,-32,15,15,17,2,-4,15,-6,-9,13,46,11,-49,-20,24,-29,-25,-9,2,-8,9,14,49,5,46,-10,30,-14,14,35,-1,17,-27,-47,-21,27,-29,64,-7,20,3,-8,0,9,30,-4,-36,42,-19,-15,6,25,-24,-22,-8,-28,27),
	(46,1,14,28,-28,-27,41,-11,17,16,49,-15,6,23,8,-33,-29,-28,14,-10,-2,55,10,-22,-6,-8,-56,13,-16,-39,-5,37,33,-10,-10,-5,-18,-32,1,-13,-26,-10,12,4,-17,-3,-14,-31,6,70,-56,-52,16,39,32,13,2,19,32,19,25,-2,-28,-2,15,14,-27,7,24,-44,3,8,8,44,8,5,-22,8,31,-11,-30,10,-3,5,-23,7,-2,-10,2,-8,-8,29,17,9,18,31,17,38,-1,32,36,-16,31,-11,-16,-7,29,39,30,-7,30,-7,-35,8,21,9,28,-10,16,22,12,-21,10,10,-6,15,-18,41),
	(37,-7,8,2,-15,-5,35,-12,59,1,21,-31,21,29,-4,-16,-58,17,-5,27,46,-14,39,4,28,29,-71,5,-2,-26,6,36,-11,11,-31,-22,13,-16,1,9,16,15,-10,10,-22,-3,-38,-47,-11,55,-26,-52,26,16,18,15,-1,30,35,12,55,7,5,-4,4,19,-20,1,-26,-10,30,15,0,34,39,-16,-26,23,-1,-4,-13,0,-24,-29,-34,9,18,-49,9,9,-25,0,-19,-19,29,-11,5,21,27,50,8,1,19,1,9,-29,46,16,-11,5,48,-31,-15,12,-9,27,1,14,-14,18,42,-30,14,-5,-34,-11,28,4),
	(2,22,43,17,-50,-37,24,-22,45,-27,-28,-35,6,27,28,-11,-38,-22,8,17,20,4,-1,-9,35,-21,-48,62,-28,-15,-1,61,-9,0,-29,-4,15,-43,9,11,18,-34,-15,14,-34,0,-18,-21,3,52,-29,-45,28,46,15,29,18,20,30,-8,71,9,27,13,20,4,-18,-17,1,-33,-4,27,8,51,59,-3,-40,23,34,-5,-13,12,-35,-11,-33,21,13,-45,-15,15,-26,22,-3,-39,21,7,2,75,45,57,5,-33,18,-21,-5,-42,39,16,8,6,55,-19,-40,-18,-6,-8,-9,-3,4,46,10,-46,30,-28,-28,0,32,44),
	(1,0,3,0,-40,-35,41,6,15,1,-11,5,-19,34,-9,-6,-10,-4,-27,-17,35,4,10,-16,0,5,-45,65,-38,-10,23,79,13,5,-13,15,18,-14,16,2,21,-20,-47,3,-24,-18,-18,-41,-18,48,-11,-11,-2,73,33,19,38,58,8,-10,45,22,14,-28,13,-4,5,-17,4,-23,10,5,17,40,43,28,-36,29,-2,-9,-13,29,-39,-26,1,-9,21,-35,4,-2,-25,18,-43,-50,-2,17,3,62,19,44,16,-62,11,0,3,-23,33,5,42,-3,37,-12,-30,18,23,0,28,2,6,59,7,-46,24,-16,4,-6,8,34),
	(37,-33,23,22,-7,13,5,-8,19,26,-6,44,-5,34,-6,-37,-43,-4,-14,-20,21,10,-19,-43,32,23,-15,39,-8,-26,22,56,15,29,-5,-12,-5,-11,6,-9,28,-15,-35,-8,1,2,-4,-44,10,30,-30,-14,19,61,34,-25,17,44,11,-11,52,21,-12,-16,-1,20,-16,3,1,-24,10,31,29,31,31,20,-25,16,-24,-33,4,-2,-52,-41,7,-13,27,-44,2,-15,-48,21,2,-34,-11,49,-13,61,11,-14,41,-16,21,22,-9,-19,5,2,22,-22,0,-30,-1,12,-2,18,36,1,16,74,-5,-8,15,-19,-11,8,-15,21),
	(41,20,30,21,-128,22,6,-10,3,-1,-38,40,-4,37,16,-1,-38,-18,17,-3,22,-13,0,-16,43,9,-17,24,-19,-11,15,14,56,41,-18,-30,24,-36,11,2,30,-26,19,-31,-10,-8,-72,-43,15,21,-21,-10,-3,62,9,-18,35,39,4,-20,72,48,-4,6,7,43,21,26,20,13,27,-14,69,-10,19,9,-15,18,-16,-18,-7,17,0,-65,-41,-24,16,-10,-18,-46,-52,15,-12,-5,31,12,-3,63,-42,-20,55,-8,-1,4,-9,-6,28,12,-5,8,6,-31,-4,10,-38,-10,36,-6,-1,70,7,-26,-4,-9,-39,15,-7,24),
	(19,15,23,19,-95,-15,12,0,27,20,-22,15,21,50,0,-13,-69,-33,22,13,30,-1,-31,-29,33,-4,-55,33,-1,-18,43,52,19,37,10,-20,13,-43,13,15,33,-51,-2,-11,-14,-1,-50,-74,18,38,16,-30,17,46,14,-17,46,58,16,-20,86,65,-32,9,-11,14,3,0,24,-15,-1,27,63,22,-2,20,-21,2,26,-44,-10,-1,-43,-29,-9,0,25,-36,24,-12,-40,-6,4,-24,14,26,-5,80,-39,5,35,-33,24,-24,-13,-26,7,31,-6,11,14,-10,-19,20,15,10,7,7,-22,57,2,-8,-7,3,-36,41,15,17),
	(22,-36,55,2,-82,-23,45,-9,18,-15,-2,-34,42,43,15,-24,-55,-24,-11,23,44,14,2,-54,13,23,-82,46,-33,-35,43,86,10,14,-17,-3,17,-78,1,-9,29,-62,21,8,-1,-15,-84,-41,4,71,-31,-24,4,68,32,24,19,55,38,-6,104,68,-3,15,23,29,3,24,4,-23,2,-13,51,29,46,35,-14,0,17,-18,-31,-4,-13,-3,-25,3,15,-19,8,-22,-68,40,22,-20,47,43,20,66,-48,0,12,-35,13,-15,-33,-43,54,40,17,26,42,0,-54,-10,-4,16,9,23,-17,46,35,-50,41,0,-34,55,18,41),
	(38,-25,39,-4,-80,-17,2,-48,-9,9,-42,10,-3,35,25,-12,-29,0,0,26,60,8,-12,-19,11,15,-31,-3,-23,-35,19,80,26,-16,-31,-27,6,-41,19,27,63,-27,-6,-16,-9,-17,-54,-15,0,7,-7,-26,22,61,42,6,4,27,19,2,76,5,-9,-21,9,3,3,6,53,18,20,13,62,18,52,35,-1,24,13,-30,-8,-12,-17,0,-15,0,25,-25,-24,-2,-31,-1,17,-49,19,0,12,15,-24,9,8,-17,22,-25,-35,-65,19,-6,-7,-1,29,-28,-24,-12,-26,30,6,32,11,60,44,-4,11,23,-36,30,25,17),
	(52,14,41,2,-90,-23,-4,-33,-22,23,-47,4,10,58,18,-4,-29,-14,-23,40,45,8,-11,-26,22,13,-54,15,-40,11,26,80,25,-19,-9,-1,19,-31,-2,-5,31,-31,0,-3,12,0,-66,-59,-14,30,26,-38,23,35,19,-15,41,24,-13,-14,41,22,-24,-25,22,15,21,6,42,-2,17,1,83,29,28,26,-25,35,-22,-44,1,9,-28,-31,-34,-9,30,3,19,-5,-48,12,7,-24,14,-2,13,35,-17,34,12,-17,-8,6,-3,-43,3,19,30,4,32,-39,-16,8,-17,-12,9,24,19,67,16,-18,-8,-7,-29,19,33,20),
	(47,-3,22,10,-40,-20,25,-37,12,-14,-35,2,-7,45,10,-23,-22,-9,13,18,22,20,-18,-34,35,3,-43,20,-23,-3,18,94,24,15,-14,14,6,-7,40,1,42,-5,-9,23,-8,0,-38,-37,16,65,-20,-34,12,83,21,-9,58,23,7,-3,43,32,-31,-1,46,-11,7,60,23,-9,14,26,27,25,37,60,-29,18,-23,-47,24,2,-72,-47,2,-11,3,-6,39,7,-40,27,25,-32,12,12,18,43,-36,10,11,-18,-2,12,-4,-15,39,28,48,-29,37,-32,3,14,-31,-1,48,-12,33,54,8,-13,-16,-9,-54,21,-5,45),
	(16,8,22,24,-54,-28,35,-49,29,4,-37,-30,23,19,15,-48,-58,-14,10,-5,44,34,-20,-33,5,15,-50,30,-23,-24,27,59,17,18,-15,-11,16,-25,26,-16,16,-28,4,8,2,-17,-58,-28,19,64,17,-28,29,45,52,-9,16,8,8,-16,41,-28,-20,20,4,0,0,31,20,-13,29,28,5,27,17,28,-8,0,7,-27,-4,-10,-23,-36,-23,-36,5,-13,16,26,-39,0,2,-43,0,13,-14,33,13,7,0,-8,1,-9,-31,-26,15,37,1,-21,46,-25,-4,12,-31,-22,39,19,26,43,5,-18,17,17,-70,33,13,25),
	(16,-1,15,25,-63,-39,6,-51,24,35,-32,-10,25,46,-4,-19,-37,-12,32,4,21,55,-8,-2,14,-15,-54,4,-5,-10,-2,61,22,19,-27,-45,24,-28,-30,22,64,-40,22,8,-28,7,-22,-48,4,39,22,-29,12,36,35,-33,-12,42,21,3,9,-9,-22,-21,17,-8,29,-29,47,34,-15,30,10,7,9,12,-18,26,-11,-35,-14,-18,-56,-56,-31,5,35,-5,5,-4,-36,-1,29,17,0,16,-33,34,6,37,18,-21,2,-19,0,-28,-2,33,7,-1,1,12,-50,8,-33,-8,44,59,-9,36,28,-22,13,26,-46,28,1,-15),
	(28,18,39,8,-71,-38,34,-15,15,8,-53,-1,37,80,-3,-39,-59,-7,22,-17,32,8,-56,-7,28,18,-22,37,-18,-9,35,47,27,4,-32,-31,28,-38,10,12,38,-55,23,0,-28,-7,-24,-25,-17,35,-31,-39,6,60,13,14,9,28,20,11,27,-8,-1,-25,-12,23,21,4,24,16,13,7,2,-5,35,39,8,23,-2,-41,-26,13,-36,-51,-12,-37,31,-8,-10,5,-36,0,29,4,25,-11,-3,64,-9,8,21,1,4,-13,-27,-56,33,26,15,-42,38,8,-9,-15,-27,24,26,-5,-10,56,29,-26,0,-12,-40,43,-2,26),
	(11,10,43,12,-66,-17,16,14,5,27,-70,-34,4,82,32,-49,-53,-8,-6,-28,48,6,-53,-7,5,3,-31,41,-40,-15,28,69,13,-22,-15,18,-6,-50,17,3,11,4,26,39,-22,2,-48,-13,-11,-15,-9,-34,9,46,29,47,8,-4,43,0,21,-16,-19,15,-35,58,12,-39,21,-3,12,-32,0,32,42,23,-11,36,30,-32,-14,17,-31,-47,-39,-14,-7,14,6,2,-15,0,3,-41,38,10,1,35,-1,36,-17,-29,-12,-40,8,-67,42,18,4,18,25,6,-16,-6,-3,-3,17,8,-11,23,18,-4,-3,-21,-33,21,13,39),
	(-10,-20,28,13,-59,-41,24,2,3,27,-31,-20,23,41,38,-7,-25,-6,-6,-27,37,33,-26,-7,19,-26,-48,35,-30,-5,11,50,13,1,5,-6,8,-49,2,7,43,20,6,-3,-36,11,-44,4,15,9,47,-22,38,27,18,-2,9,3,20,-16,46,-7,-10,-5,0,33,-9,9,-6,57,9,-19,-41,16,5,16,-40,17,4,-8,-7,-22,-48,-5,-29,-14,14,8,-4,-10,13,-6,24,-10,44,23,-6,35,-19,47,-1,-15,2,-23,-5,-40,16,7,-5,13,11,-3,-45,16,-15,-18,30,22,-4,26,-7,0,0,15,3,18,1,6),
	(27,23,-5,-6,-63,-18,18,-28,-8,18,2,-32,-2,34,29,-14,-4,-2,-19,-9,2,5,24,2,-9,-4,-34,0,11,0,-18,17,22,30,-25,-20,-5,-14,2,-4,15,-1,39,19,-4,-19,-24,-29,-5,23,13,-35,9,35,1,18,17,16,52,-7,11,-2,1,-2,-17,43,-29,37,-11,2,-9,-8,-50,21,28,0,-28,10,12,-26,-18,0,20,-7,-28,-22,8,-21,25,2,-16,31,-28,-23,41,1,-26,26,-23,39,33,-11,1,-38,-11,-52,42,-17,-7,-4,43,1,-9,20,1,-2,-3,-16,20,12,-7,-9,2,25,-22,4,-6,36),
	(5,11,-11,-4,-8,10,37,-14,16,2,17,-37,18,34,15,-8,-43,-22,-20,15,4,20,30,20,-28,36,-36,0,27,15,-25,7,-18,-12,8,18,-6,-12,-7,13,-11,16,38,-17,-15,19,-18,-41,-19,26,-45,-21,-31,24,16,7,-4,-5,42,9,0,-11,13,18,-8,28,-2,16,-37,-21,44,0,5,15,27,41,-32,-10,23,-19,0,18,18,-19,-17,34,-15,-20,6,-20,-19,26,-36,3,25,-14,8,7,1,-7,4,-22,-19,-27,-2,-36,34,19,6,16,23,15,-15,-11,-15,-5,20,0,-13,14,10,-11,13,-21,-6,8,6,8),
	(9,-5,-9,-10,-1,-3,-6,16,-9,0,-9,15,2,0,-1,21,-18,17,-2,18,9,0,10,14,-4,-14,7,-14,-11,-8,0,4,15,5,16,0,14,-12,-11,0,10,0,9,-3,-7,-14,-13,16,0,-4,-9,5,17,-13,11,19,0,1,-6,-6,-3,10,5,-2,-8,11,11,-11,-2,27,-3,19,-18,0,4,-3,-11,-10,-11,9,-10,-13,7,23,-7,12,-10,-1,1,-6,2,13,1,-22,5,-5,-2,-5,20,17,9,-8,-19,17,-12,16,9,-8,9,4,7,6,-14,20,-12,-20,-13,11,2,15,-11,1,-19,10,9,17,21,-22),
	(-4,-10,6,11,1,4,15,-12,1,-17,0,-18,11,5,-19,0,-11,-11,10,2,16,-18,-12,10,19,6,-16,17,-4,2,16,-1,-9,15,-9,-18,12,17,11,-13,15,-15,6,5,-7,-5,6,-2,7,9,-19,-15,-18,7,6,7,17,1,-2,-16,-6,6,2,-7,-1,7,-5,7,16,17,11,8,14,12,-16,-8,-6,15,-9,20,16,-9,-20,-20,-17,14,9,18,0,20,-12,19,-7,-18,-19,-11,18,-18,-2,14,4,10,0,8,-15,5,4,-14,6,-10,0,-3,-11,0,9,-12,12,4,8,-9,9,-10,-16,12,-19,-11,-4,16),
	(17,10,7,-19,12,-3,11,19,14,-16,12,-11,-13,12,10,-4,-6,18,-12,12,-9,-8,19,-16,14,-5,-10,19,20,-7,-9,16,-11,-2,-9,20,8,16,18,16,16,-16,-5,-4,-18,-6,-18,-1,2,-13,15,12,3,17,-6,3,10,15,-3,6,-15,-14,9,-5,7,-19,17,-7,15,12,12,-4,2,11,17,0,-1,-18,11,-14,-16,-4,-3,-5,-16,-12,-13,0,19,9,12,5,13,18,-1,17,4,0,-15,17,12,-15,8,-17,-11,-17,0,10,-16,-16,13,16,-5,-2,0,10,-15,3,2,-18,18,-18,-11,-1,-19,-2,20,-7),
	(-9,-13,-3,-7,-17,-1,-10,-11,7,15,-10,-17,5,18,18,-5,-15,17,3,-8,-12,-17,-7,-20,-14,13,2,-13,-15,11,-16,0,-5,-4,12,12,16,-12,12,-13,9,-8,7,-7,-6,-17,16,-17,-19,-16,-6,-18,-6,-6,-1,-9,16,-6,-10,0,6,17,-1,4,-9,12,-2,9,-3,17,-9,10,11,18,9,-6,-11,-2,18,-15,-11,-4,13,-19,4,10,17,-13,4,-15,12,-15,9,-16,-10,11,17,2,5,-20,15,18,1,-12,6,19,-11,-5,1,-5,-16,14,4,-20,-15,0,17,-9,4,5,19,10,-3,-6,-17,-2,-18,1),
	(10,0,10,-10,0,0,18,12,-18,-5,16,16,5,15,4,14,-19,-15,13,11,15,3,15,-9,0,-1,-15,5,18,16,8,-12,9,14,-1,14,2,-10,0,9,-7,-16,-9,-11,1,-19,6,-7,15,-2,-1,-5,-7,9,-2,10,3,6,12,-2,-12,-4,12,19,-20,11,-13,3,-12,8,-3,20,-12,5,1,-9,4,5,18,0,-2,8,12,19,-13,13,-20,-8,-5,13,6,18,-12,-11,-13,-14,10,5,9,20,-18,14,16,8,0,16,-5,13,-8,-4,20,0,3,13,-7,3,-17,-2,5,-16,-9,11,-8,13,6,-20,-9,19),
	(-7,10,14,12,17,3,1,-6,19,-9,19,9,7,19,18,17,-12,-3,-15,-14,-9,17,-20,5,4,-20,-19,6,-16,16,18,-1,4,1,-9,-7,-10,8,-15,-17,-12,2,9,-19,2,0,-18,11,-9,15,-17,17,1,11,-17,10,13,4,-2,7,-15,-12,-9,5,-13,-6,20,-5,-20,-7,-20,-11,-15,0,-12,2,-14,-8,-11,1,-19,7,17,13,2,0,-5,-17,0,-3,10,13,-13,12,9,3,5,11,-19,-1,-16,12,-2,-1,-8,16,11,-16,0,-5,9,17,-20,-19,13,2,-8,-15,-13,-18,-4,13,15,6,-14,6,-12,-2),
	(-2,-1,1,-10,7,-17,6,0,-14,6,9,-13,-4,10,-4,11,3,-8,-13,-1,14,6,-5,-1,7,-14,-20,11,0,5,2,7,-13,-16,-11,-17,4,8,-2,-5,-9,-4,6,2,16,-8,-2,-17,-11,7,-6,2,-5,-4,-1,-14,5,10,-15,0,15,-6,-2,10,-17,-5,-9,3,-4,-16,18,-4,12,3,5,4,10,17,18,9,17,19,-17,-6,17,-18,20,-2,-12,-14,17,-3,11,11,-15,20,-14,-1,-11,9,-14,19,-9,1,-11,20,16,-10,-19,17,-11,15,-10,-7,18,-8,3,-12,-16,-11,15,-13,16,-16,13,7,14,-15),
	(13,15,-13,5,6,-9,-30,13,-11,8,17,-7,1,-28,-15,-18,-4,0,7,-11,8,13,2,-9,-12,-3,21,-31,3,-13,-5,12,-8,-13,32,17,11,26,3,24,15,-5,2,-3,-15,-16,2,-8,20,17,12,11,25,-20,0,-2,16,8,-1,15,-25,11,-7,-10,-9,17,-12,-11,10,2,-3,14,-3,-6,-17,8,-22,-32,8,15,1,-22,0,31,0,10,-13,12,-5,-4,0,-8,8,-13,-27,0,-2,-28,-9,17,-10,0,-23,-21,0,6,-27,14,-19,-15,-23,6,-7,28,-7,-29,-4,6,-24,2,22,10,-6,10,31,-17,-9,-33),
	(-17,-7,4,-13,-5,2,-26,12,-15,0,27,-11,-3,-21,22,-11,-12,17,26,17,-5,20,16,-14,0,-16,-6,-29,20,-16,-12,14,-5,18,20,-12,20,32,-4,3,-1,0,17,-9,-22,-12,19,-17,18,-6,5,-5,-4,-1,-14,13,-16,-7,0,4,-1,8,16,1,7,-12,-27,-11,17,34,-18,6,-6,8,9,-31,-13,-6,5,17,11,-24,-18,17,11,10,-1,-10,11,11,-8,-2,13,6,0,-20,-3,-11,-16,30,-16,-20,4,-31,9,-4,-30,21,-36,-8,-22,-5,-26,21,0,2,-25,3,-20,5,-2,11,15,45,23,-10,-4,-26),
	(6,-18,18,-35,-5,-16,8,-14,1,-3,62,-13,26,34,-9,21,-7,37,12,-4,6,34,-19,-9,3,8,-23,-5,-6,-7,5,25,-3,8,22,-26,-4,-16,-23,-17,25,17,31,4,-31,-18,17,9,-7,2,-17,-13,3,16,6,9,3,41,11,-19,13,6,20,-21,-3,29,-3,11,16,-2,8,14,-9,6,-3,-10,-25,-17,-7,-29,-26,-10,-32,-4,-23,-14,-13,11,-13,-4,-6,3,41,-5,20,3,-1,12,7,36,12,5,28,-33,-8,-13,19,7,-22,10,34,-17,-26,-14,0,8,2,27,-5,14,7,-5,-4,38,-20,-3,7,11),
	(41,0,24,-23,4,-7,29,-17,0,-14,57,3,6,41,14,-6,-27,1,10,7,12,18,4,-14,33,11,-9,18,-12,6,-4,25,20,-2,-15,7,14,-8,-4,-16,8,-7,-3,6,-20,-14,-11,-11,-2,30,-18,-4,-12,-5,15,0,17,38,-2,8,14,18,13,7,-38,37,8,-7,22,11,-5,15,14,8,-5,18,6,11,1,-1,11,4,-25,16,2,-5,-12,-20,-14,-20,-8,1,10,27,26,-11,-2,12,0,-6,25,-32,13,11,-31,-17,2,7,-23,-17,23,0,-23,5,12,21,-18,22,-7,1,15,-15,2,7,-6,-12,16,-4),
	(20,-10,-6,-1,-29,-15,35,-20,2,-27,66,2,-4,34,20,3,-40,-12,21,-6,25,20,-21,9,35,25,-26,28,-27,22,-13,3,9,0,16,6,7,-24,1,-24,21,7,0,28,-24,1,25,-24,-21,20,-36,-32,24,-14,2,-8,22,19,34,-12,20,4,4,2,-5,18,26,-7,19,13,-14,-4,40,24,-22,14,-20,-10,-15,3,1,-7,0,-11,-7,3,3,-25,-3,-13,-32,14,15,5,27,-9,0,19,-7,-11,10,4,19,-17,-19,-37,3,18,-22,-21,20,-18,-9,7,-32,17,-7,5,12,0,-9,-2,7,13,-20,0,23,-9),
	(-5,-21,-7,-1,-3,-24,29,0,-5,-5,56,1,21,54,-8,19,-14,0,3,-8,40,37,-6,-9,9,-3,-12,-8,0,-14,-15,21,12,13,18,-3,9,-15,10,-7,35,16,6,21,-10,-8,12,-11,-9,20,-31,-16,13,-9,1,16,18,6,20,11,8,17,-3,12,-7,33,9,-21,42,16,4,-4,11,19,-14,-4,-28,3,19,0,-11,9,3,8,-23,24,-5,-27,-20,-18,-11,-18,54,9,22,-4,-9,-3,-1,-1,18,-45,14,-11,-8,-39,-7,-2,-24,3,31,-16,-21,0,-3,14,4,2,-18,3,0,-11,15,44,-11,-10,18,10),
	(3,-1,29,19,-9,-22,33,-33,36,-22,3,-19,16,50,34,5,-42,29,26,12,33,16,27,-22,23,-22,-11,32,-17,3,-4,35,-24,0,-9,-40,12,-11,-26,8,28,21,44,22,-35,12,51,-27,10,33,-60,-38,25,-3,5,-1,-12,23,12,16,19,1,-26,-8,23,49,9,-38,26,11,-2,44,45,16,0,-8,-29,6,31,-13,-28,-19,-33,49,-21,5,33,6,13,-6,-13,-2,31,-11,7,-5,-17,13,5,35,10,-21,7,-37,38,-44,0,15,-25,17,29,-7,-28,17,-24,41,-26,28,-36,-2,14,-6,53,12,11,-34,52,-9),
	(0,-30,26,6,-45,-12,31,-8,4,-27,23,-17,24,62,18,-9,-35,16,3,5,46,28,44,-1,30,13,-46,14,0,14,-3,34,11,-4,18,-8,17,-19,9,16,21,22,23,-9,9,-5,1,-23,3,1,-55,7,0,24,0,14,21,3,13,-20,15,-16,-1,-11,37,28,25,6,13,-1,0,8,28,-3,12,19,7,7,5,-3,-9,0,-25,48,-5,-16,8,5,17,14,-33,-16,54,-18,21,-6,-2,19,17,-5,-1,7,15,-15,-8,-52,3,-1,0,-6,-5,3,-10,-17,-4,32,-19,21,11,12,8,17,14,20,-22,-4,22,-14),
	(3,-51,17,4,-8,-15,2,-40,-12,-9,-5,-16,15,27,9,28,-30,1,6,-17,21,14,-7,7,25,-3,-3,29,-12,15,3,22,16,-8,-13,-24,6,-1,-10,5,38,-23,35,5,-9,-28,-27,-15,20,9,-14,-15,24,30,-4,18,17,-5,11,-4,45,-12,-17,19,11,46,7,-16,1,7,-19,9,43,0,8,-10,0,-13,-1,-22,15,4,-22,2,-23,21,9,-21,-5,0,-17,-12,15,-5,19,-14,-18,27,-10,-6,1,0,18,-21,10,-35,8,18,-8,23,30,-20,2,-16,8,18,-18,-5,6,20,9,16,-5,38,10,0,26,19),
	(0,-41,11,-45,-48,-25,37,-34,30,4,33,-26,15,49,13,14,-49,3,34,34,17,57,44,-27,14,-25,-15,19,6,7,-7,31,-11,-15,27,-9,40,-6,-12,28,59,-12,63,8,-26,27,14,-33,20,36,-23,-21,30,22,2,10,-35,40,14,1,12,-11,-17,-3,-34,21,0,1,-1,43,-33,43,-11,23,-6,-27,-20,7,8,-17,-30,-40,-19,2,-15,37,30,-7,-10,3,-8,-2,65,-4,34,0,0,10,10,38,10,-52,-14,-2,30,-49,-11,28,-45,17,23,-11,-47,16,11,-17,-31,34,-23,35,12,6,28,46,11,-7,33,-11),
	(33,-19,16,-2,-61,-28,26,-38,32,-11,19,-47,12,77,20,-6,-53,25,3,17,64,80,24,-12,44,12,-44,-1,-9,-19,26,68,-4,8,6,-9,0,-45,5,-27,18,-1,43,59,-24,-37,-10,-43,3,33,-64,-50,35,56,5,12,19,46,63,12,35,-15,7,5,52,46,46,-2,4,-31,23,13,41,48,13,12,-26,35,33,-24,-25,-18,-26,-17,-5,-17,-13,-52,-6,-37,-28,-6,76,-15,41,49,28,56,-5,36,-10,-10,23,-8,7,-54,28,44,-18,0,62,-67,-32,-11,-22,7,-1,15,-18,56,6,-1,29,14,-6,12,37,12),
	(28,-24,27,0,-55,20,-4,-16,21,-10,10,-47,5,43,0,-4,-38,26,21,9,23,13,45,-9,30,-2,-31,-9,-22,-26,20,40,-2,-10,-14,20,6,-31,19,-11,-9,6,7,44,5,-15,22,-1,-2,25,-9,-27,20,24,2,21,3,-6,13,-9,50,14,-23,5,17,45,16,11,34,-17,16,-8,37,31,15,38,-4,18,0,-13,13,-8,-3,0,-27,-16,7,-30,20,13,-51,29,5,-7,22,34,23,41,-5,54,-6,-7,5,4,0,-21,24,12,28,-9,28,-62,5,-27,-6,15,19,0,21,7,7,-21,36,-19,-31,7,31,22),
	(35,-24,12,23,-27,-2,34,-66,17,-7,32,-45,7,16,47,-12,-27,41,28,0,16,3,-4,-12,39,0,-40,-18,4,31,1,30,-16,-1,-10,2,23,-50,-3,5,38,20,15,13,-7,7,25,-24,3,52,-19,-35,24,36,7,0,-12,15,41,7,38,-7,-22,-26,42,27,-2,-1,5,10,-11,-1,11,23,8,16,-9,-18,22,-1,-16,-33,-17,40,-49,12,18,-36,15,19,-4,-5,32,1,29,1,31,31,1,36,-1,-2,-23,-21,26,-47,-9,44,-30,8,7,-29,-19,15,19,8,-11,18,3,24,31,-20,29,12,-22,11,46,-11),
	(32,-6,18,-2,-25,-33,38,-43,11,6,-17,-50,4,0,41,20,-13,12,6,13,28,68,34,-14,18,-46,-10,0,0,-7,-24,47,-13,-12,-15,-15,43,-23,-14,28,46,-9,53,-16,-14,-16,-21,-30,10,31,-17,-41,20,6,29,0,-8,29,34,-18,0,-15,14,-16,0,34,18,-19,37,13,-30,19,-20,37,2,0,-8,0,31,0,-35,-10,-25,-17,-42,42,39,-17,-3,7,15,-20,34,8,28,-12,-9,9,1,21,-21,-17,-11,-19,0,-18,-2,30,-3,26,27,-22,-52,26,18,15,-21,10,-26,28,8,-5,40,63,4,-15,0,2),
	(20,11,36,15,-52,-8,24,-68,1,0,-43,-30,17,35,36,-12,-3,-15,-12,21,18,17,9,6,33,-6,-21,0,-1,18,21,30,1,-14,0,-16,20,-3,0,-8,-7,-17,43,36,11,0,-4,-35,14,25,0,0,4,38,-10,13,-12,34,43,15,29,-17,10,-7,21,42,11,-20,-13,-20,19,-22,-5,29,26,-4,5,18,13,3,-2,13,2,-27,-34,33,-15,-19,-4,-39,0,-10,39,-8,58,-13,-33,7,-8,8,1,4,-9,12,15,-64,9,0,-1,30,20,1,-37,3,-19,-2,14,-2,16,1,3,-8,30,29,-17,2,0,-6),
	(0,14,23,-5,-41,0,47,-50,-3,-5,-24,-26,2,1,4,-33,-15,-23,12,15,10,5,-8,0,39,-12,-30,21,-23,-15,24,42,-11,-8,-2,4,8,-10,24,-16,21,-13,0,19,-23,-10,-30,-29,-24,24,-16,-13,2,10,7,21,-1,8,49,14,11,-13,12,16,10,9,6,-11,-28,-18,-7,-8,-19,31,3,-10,5,8,13,-2,17,16,-10,-34,-42,11,-7,-10,12,-28,-15,22,48,18,51,-8,-22,25,-10,-2,-8,-26,-16,-19,19,-22,34,-2,17,25,52,7,-34,-29,-19,-1,2,13,-10,1,-2,-6,20,19,-28,24,-2,24),
	(-10,5,-7,8,9,2,20,-19,-21,10,-31,-16,31,22,6,0,0,-22,-17,0,21,27,26,-14,-9,-13,13,12,-2,6,-24,0,13,7,-15,0,29,-7,6,4,-1,4,-12,31,-2,5,-23,-9,19,-3,-18,-5,-8,15,20,9,-18,11,24,-6,-9,13,7,8,-11,2,16,-7,-28,26,-19,3,-27,26,-7,-1,-13,19,19,15,-11,4,3,9,-17,-10,-8,4,1,3,-11,-32,-22,3,19,8,-21,-13,16,-8,-23,1,12,-19,0,-1,5,-16,-15,7,-2,0,-7,-1,-3,-1,8,-9,5,-6,0,-2,33,11,-4,-17,-1,-18),
	(5,-24,11,25,6,-6,29,-19,-13,22,-51,-45,26,6,37,2,6,-3,-10,-12,19,38,0,-6,-25,-1,-34,-5,-6,-13,-19,36,-14,-47,0,-13,16,-25,-39,-2,24,16,34,14,-24,0,-27,-27,4,-9,25,-24,38,-14,-25,45,-1,14,45,9,-13,-17,-17,-18,-15,16,18,-8,25,31,-35,-3,-13,18,-24,-44,-32,-11,28,-9,-27,-13,-22,6,0,38,23,-11,-21,-17,24,-41,-43,1,17,0,-4,-13,-6,38,-6,-39,16,-9,17,-29,23,5,15,38,31,-26,-28,26,-10,16,-4,14,-16,3,-12,-22,-2,18,38,-9,7,-26),
	(-16,-20,-5,28,-14,-4,20,20,9,42,-39,-38,9,13,24,-22,-16,5,-37,14,17,45,-32,-3,-33,-25,1,10,13,-8,-10,40,14,-42,19,4,30,-26,-6,10,26,31,22,56,-22,14,-44,-20,14,-5,48,-16,41,8,-31,13,-29,4,28,8,-15,6,-22,-11,-13,12,19,-26,18,14,-24,-25,-26,45,-18,-47,-9,10,36,30,-1,-38,-7,-9,7,36,6,-18,-16,12,24,-20,-13,-16,16,17,-11,-5,17,29,-32,-30,8,0,30,-3,-14,-16,-16,51,35,-1,-2,26,24,7,-6,3,3,-22,-13,-10,4,33,12,-32,-22,2),
	(10,-6,27,12,25,-33,-5,-12,-1,31,7,-28,5,25,37,15,6,37,9,-8,12,44,17,15,-38,-37,2,18,7,16,-21,-5,-10,15,24,-9,33,-3,4,34,28,5,6,7,-35,-19,-15,-3,37,24,40,2,20,-28,-14,34,-5,-7,-4,0,-4,6,-16,-30,19,6,0,12,9,31,-37,19,8,8,-16,-21,-38,-15,4,18,-18,-34,-21,0,1,25,19,-11,6,-1,-2,-4,28,-6,6,-12,12,17,-16,32,-33,-6,17,-15,-5,-18,-18,1,-12,11,29,-16,-8,5,33,-26,17,-7,6,0,17,-32,10,14,-6,-4,22,-34),
	(-4,8,18,0,0,-13,-14,-17,0,-4,12,20,-12,-10,14,-14,7,-11,3,-8,-7,-16,12,-6,-9,-9,-11,-7,12,-16,17,-7,-12,-12,7,-13,12,11,-1,16,-19,1,-16,15,-13,4,1,-11,-1,12,13,-8,-16,-11,1,4,20,14,0,4,0,11,2,17,12,-13,-14,10,-14,2,-8,0,-7,-8,-9,-18,0,16,-3,3,20,-6,-17,-6,-18,16,-19,13,0,-9,-17,12,15,13,-13,-7,13,-2,13,11,17,9,-17,0,0,7,3,-5,2,-12,16,-11,7,5,-1,-16,-4,12,6,12,-9,17,10,1,16,-19,18,20),
	(6,-19,5,-16,16,-10,0,-4,1,-13,5,-1,0,1,-15,3,-10,-2,-8,1,-16,11,15,6,-4,-18,12,18,11,-1,-13,7,-12,-15,-14,-14,-2,7,-7,-8,12,0,-10,-19,-3,14,-2,-6,0,2,-11,-3,17,-17,-19,4,13,5,6,-11,10,15,-8,19,11,0,-10,-16,-1,-1,8,-16,4,8,-1,-3,-18,18,7,3,-16,0,0,1,9,-19,-20,-11,0,-19,1,7,3,-7,20,-8,3,3,-17,-7,-10,-3,5,6,-10,19,18,-14,-13,13,-18,8,0,-18,-11,2,-3,18,-2,2,-8,-20,-9,-3,-8,0,-3,-11),
	(19,13,-1,-16,-17,3,-15,11,8,16,7,-5,-10,-18,14,11,15,15,-12,19,4,7,-18,-1,-3,17,-6,-8,-8,3,11,14,9,6,-20,8,-9,-8,-10,-7,-4,-3,-12,-2,14,17,0,5,-1,-8,2,10,2,17,-6,-1,1,-19,-13,14,10,18,0,3,11,-12,6,5,-18,-9,-11,17,-20,16,-4,14,4,19,-19,0,8,-20,11,19,4,10,-12,-6,17,-17,-8,-16,7,14,-1,19,11,-11,-11,-14,-12,-12,20,-1,-12,17,18,-17,-7,-2,8,-7,3,2,-3,-2,-17,-18,1,11,9,3,12,-14,20,-6,10,-13),
	(11,-4,-14,-6,18,-2,1,-18,3,-2,-15,4,-3,14,18,15,-17,6,-7,18,-5,-8,10,-2,1,-20,-1,0,14,-15,8,-4,-18,16,-20,-18,16,15,-13,-14,0,1,-18,-9,-10,-9,11,-10,17,12,1,-16,8,-15,-3,13,2,14,-5,6,15,-8,10,-20,17,-15,8,10,-12,11,0,17,-3,-13,-13,13,18,1,11,-6,-14,-16,19,-2,-19,5,-12,4,13,-8,20,7,-19,0,-14,4,-12,16,-18,-16,-5,-16,10,3,-11,12,-16,-14,-4,14,-2,-1,1,-13,-4,-17,13,6,-10,-16,18,-1,-10,-1,2,7,20,4));


	constant weights_2 : weight_2 := ((-144,-17,42,-126,-37,65,89,-113,-10,71),
	(82,-52,-185,15,59,21,73,-2,-129,80),
	(-82,-28,-52,-4,61,81,-163,56,-51,64),
	(-2,38,58,6,-107,-50,-43,-39,35,-8),
	(-43,101,-136,-105,157,-33,42,-38,-52,-128),
	(-59,39,43,-18,47,-20,59,-90,17,-19),
	(50,-70,53,-53,-2,-50,22,27,48,52),
	(1,-10,1,46,6,-2,-33,-90,90,-23),
	(-80,20,32,26,5,-52,-70,29,42,18),
	(62,-7,-14,73,-6,-37,24,96,-103,-97),
	(-33,84,126,35,-39,8,-8,-1,11,-164),
	(66,-42,-67,20,-50,86,32,-60,48,-55),
	(-47,58,55,11,-98,0,-88,38,-4,35),
	(-4,97,-63,-36,-54,65,-63,43,-148,97),
	(-71,-50,9,-105,49,-116,86,75,-27,30),
	(28,-29,62,-24,-101,-1,10,-7,-40,-107),
	(13,2,47,44,60,-54,23,-23,-42,-107),
	(5,34,42,-22,-107,0,-42,17,44,-53),
	(-110,-6,17,0,-68,-19,-33,55,37,-89),
	(18,-52,48,42,27,3,-53,31,-51,-69),
	(-9,26,14,-45,-134,65,-175,56,-8,32),
	(67,44,3,-92,4,-22,-62,165,-16,-9),
	(78,109,-1,-16,114,-93,-4,44,-108,-14),
	(42,33,-81,-138,62,-39,-33,6,63,5),
	(54,-65,-28,-55,-19,51,-14,12,14,23),
	(-55,20,44,16,-8,-6,19,-47,40,7),
	(-69,72,-24,-34,89,37,-72,-36,4,-116),
	(22,-18,60,39,-132,-40,-29,14,-14,55),
	(-101,50,31,47,55,-116,48,56,1,-51),
	(58,30,-80,16,-94,90,77,-18,-76,-119),
	(-64,29,50,-4,-1,57,-11,-37,23,41),
	(-43,24,-52,54,-50,-6,87,6,-40,20),
	(43,-72,45,52,6,42,-7,5,27,35),
	(45,80,-89,-33,-72,90,97,-40,4,38),
	(-38,40,51,-41,35,42,23,41,44,-19),
	(-127,50,-40,50,44,-55,-63,-101,63,15),
	(-3,-77,10,-40,-8,53,-3,55,-21,5),
	(-69,57,29,48,61,53,-55,-8,39,-53),
	(-86,46,-123,16,64,46,5,-38,-34,40),
	(-31,-35,-34,57,37,56,-42,46,-34,-25),
	(35,90,-51,5,-78,76,-57,30,-87,-24),
	(-127,52,-19,-80,26,55,41,60,34,-51),
	(140,26,88,-25,-69,-191,70,52,-11,16),
	(69,52,55,-29,-11,-114,60,-8,6,23),
	(-38,-73,-6,21,49,16,-5,-71,36,7),
	(-44,75,-31,25,80,-27,31,62,-105,-27),
	(35,17,31,12,-50,-33,63,60,36,-176),
	(-87,94,48,-103,6,49,54,-38,66,-122),
	(0,-79,-56,30,28,42,-28,43,34,-23),
	(-16,-50,-59,20,-10,-70,41,22,8,9),
	(48,18,21,25,-46,-51,-33,-15,103,-139),
	(43,-28,42,30,54,32,-23,-40,37,-15),
	(37,-48,-37,-78,-59,-10,-20,45,29,-29),
	(-44,44,-2,44,-56,47,-97,19,7,73),
	(-49,33,33,63,16,41,-151,55,-30,44),
	(-59,24,52,4,64,-32,-57,46,31,51),
	(-19,-5,-123,19,25,68,15,3,50,65),
	(29,-75,0,43,-69,-44,-76,28,-28,2),
	(49,-74,-51,-31,-12,-53,-49,20,-1,16),
	(0,42,16,-32,-6,-50,29,43,38,-46),
	(17,-36,-42,37,-75,14,-16,-5,20,28),
	(-16,60,110,94,-107,45,-129,99,-133,-69),
	(38,32,69,17,8,-72,-89,87,-4,-56),
	(16,66,-1,-21,45,-66,14,-55,31,14),
	(3,63,-102,-105,58,-109,-98,-35,-97,119),
	(51,-106,-34,-56,30,37,7,41,32,45),
	(23,-42,-158,-46,-86,100,-35,-39,10,-6),
	(3,-23,0,10,-36,0,66,-103,26,-29),
	(-81,-136,11,171,-117,51,-131,81,-100,-48),
	(25,5,-5,-47,52,70,-9,83,-8,-127),
	(-43,39,16,36,-33,-37,14,-71,45,8),
	(-20,49,12,41,-103,4,-47,26,10,-49),
	(10,-13,-63,70,-129,120,62,-28,-46,26),
	(74,16,32,57,-12,-119,-112,58,-12,47),
	(-140,36,-48,28,-48,13,11,-30,12,12),
	(-66,-93,78,81,-33,36,23,-77,-108,53),
	(-45,-66,42,-55,40,39,4,-29,35,14),
	(18,-34,61,56,-115,5,-65,-13,-21,57),
	(-10,-67,7,-46,54,-64,14,65,-6,33),
	(17,-50,34,16,52,-52,0,19,20,-42),
	(21,55,-69,-57,58,32,23,-69,8,14),
	(8,-72,14,25,22,30,-1,-41,27,46),
	(14,38,118,-13,71,-65,31,-66,-116,19),
	(-31,100,-86,6,66,-64,-22,93,-137,-169),
	(32,68,12,40,-59,5,-43,-84,21,-36),
	(68,-5,10,-25,48,-6,19,41,-112,27),
	(-118,-17,23,-8,41,106,-172,47,-178,-2),
	(-77,10,7,67,11,69,20,-43,-41,-44),
	(8,-50,-34,28,27,-22,83,-31,24,27),
	(-49,78,-6,92,1,-165,-10,47,-50,-74),
	(-18,111,-38,-110,63,5,61,23,-86,-49),
	(41,-82,-38,27,-74,-1,8,-75,34,28),
	(-3,-189,-40,-105,-119,161,103,7,17,7),
	(58,120,33,-20,0,-93,25,-80,-30,-17),
	(26,-89,-14,-67,-8,-74,-108,24,42,64),
	(-47,-160,-126,15,-76,29,-18,-74,-21,98),
	(-95,-8,14,124,-70,-47,-107,-72,-2,83),
	(-30,-122,27,25,2,25,32,12,24,35),
	(-56,23,-111,20,16,97,67,-48,-101,-191),
	(-34,-35,-47,66,72,-185,-23,119,1,45),
	(-13,-55,69,-38,21,29,50,-116,20,35),
	(-28,-56,-67,-118,36,37,28,-97,98,-38),
	(62,-51,-4,56,-97,1,40,-72,28,50),
	(-9,33,8,4,-33,-7,-27,-94,55,-36),
	(-20,43,-2,-109,-13,23,-35,36,54,-66),
	(44,3,50,0,-20,-44,8,-58,60,-57),
	(-33,-4,-59,-16,29,-45,-105,4,30,63),
	(-26,-96,-20,-5,-33,-138,97,40,43,18),
	(-25,51,-108,64,71,-72,-82,0,-81,60),
	(49,-53,16,-73,38,-13,12,27,-14,20),
	(-15,0,-9,-6,12,-18,-70,22,43,35),
	(67,73,74,-74,49,25,-36,-75,-136,84),
	(-29,-41,-11,17,9,2,60,-69,47,-40),
	(-33,-34,-39,55,8,-5,-46,11,40,-35),
	(-106,-30,10,72,39,-40,-114,26,47,0),
	(69,-19,66,22,-88,-95,27,-50,-10,75),
	(14,-40,18,47,-18,7,52,-12,30,12),
	(29,32,34,41,-81,65,-130,19,-67,-56),
	(-10,4,-116,-6,62,45,-108,-48,0,55),
	(5,-2,4,61,-105,38,-100,0,-14,5),
	(-33,-51,28,-22,-88,68,20,34,-57,-115),
	(31,24,42,-92,37,42,20,-15,11,-10),
	(-21,5,73,-124,-23,-70,18,22,-34,36),
	(-146,131,168,-63,-12,-91,42,112,43,-149),
	(60,9,92,-24,40,-8,58,44,-139,-43),
	(47,-13,-21,-39,-115,43,82,-50,6,40),
	(0,-64,44,-46,-131,14,24,45,-10,-70),
	(-34,9,-56,33,37,6,-82,0,-6,62));
	
	constant bias_1: intermediate_output := (34,-22,43,-13,19,28,0,7,-5,6,12,-5,13,28,27,24,0,8,-4,5,32,15,-1,-3,19,11,34,-12,3,11,33,0,-11,-2,29,-4,28,19,18,15,18,30,11,4,10,5,-22,28,12,-27,-12,11,1,4,7,30,10,-22,-19,-3,-18,14,-5,-14,17,18,24,-19,0,31,-11,-7,9,-8,0,11,34,-19,11,-8,7,-9,26,14,-5,5,30,18,-15,-4,19,-42,12,-8,-1,1,0,9,-2,-6,17,4,-35,-5,19,-10,0,1,0,19,0,9,-1,-14,9,-29,-31,7,15,-8,19,40,21,20,11,-16,21,7);
	constant bias_2: final_output := (-33,6,20,-23,13,30,-14,6,-4,-12);

	constant image_0: image := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,44,105,114,254,210,93,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,22,60,148,229,253,253,253,253,248,99,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,188,253,253,254,253,253,253,249,149,112,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,15,191,253,253,253,254,253,253,253,178,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,163,253,253,253,253,254,253,253,253,245,207,36,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,72,232,253,253,248,134,74,204,253,253,253,253,134,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,224,253,253,253,128,0,0,29,206,253,253,253,253,94,0,0,0,0,0,0,0,0,0,0,0,0,6,161,251,253,253,168,4,0,0,0,23,253,253,253,253,248,56,0,0,0,0,0,0,0,0,0,0,0,130,253,253,253,253,49,0,0,0,0,4,129,248,253,253,253,59,0,0,0,0,0,0,0,0,0,0,0,164,253,253,253,173,6,0,0,0,0,0,0,224,253,253,253,59,0,0,0,0,0,0,0,0,0,0,0,165,254,254,242,71,0,0,0,0,0,0,0,226,254,254,256,59,0,0,0,0,0,0,0,0,0,0,50,238,253,253,223,0,0,0,0,0,0,0,0,224,253,253,232,45,0,0,0,0,0,0,0,0,0,0,60,253,253,253,223,0,0,0,0,0,0,1,87,243,253,253,163,0,0,0,0,0,0,0,0,0,0,0,60,253,253,253,237,57,0,0,0,0,0,15,253,253,253,253,93,0,0,0,0,0,0,0,0,0,0,0,43,227,253,253,253,238,57,0,0,0,0,148,253,253,253,173,6,0,0,0,0,0,0,0,0,0,0,0,0,147,253,253,253,253,227,60,0,18,61,227,253,253,249,223,12,0,0,0,0,0,0,0,0,0,0,0,0,15,253,253,253,253,253,232,134,205,233,253,253,253,143,0,0,0,0,0,0,0,0,0,0,0,0,0,0,10,163,243,253,253,253,253,253,256,253,253,210,120,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,97,120,232,253,253,253,254,242,199,31,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,56,104,104,104,256,105,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

end package;