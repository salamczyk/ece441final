library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package project_package is
	type weight_1 is array (0 to 783, 0 to 127) of signed(17 downto 0);   
	type weight_2 is array (0 to 127, 0 to 9) of signed(17 downto 0);	
	
	type intermediate_output is array (0 to 127) of signed(17 downto 0);
	type final_output is array (0 to 9) of signed(17 downto 0);	  
	
	type image is array(0 to 783) of signed(17 downto 0);
	
	constant weights_1	: weight_1 := (("000000000000010001","000000000000000110","111111111111110100","111111111111111001","111111111111101110","000000000000000000","000000000000000000","111111111111111011","000000000000000011","111111111111110001","000000000000001001","111111111111111100","000000000000000110","111111111111101101","111111111111110000","111111111111110110","111111111111110000","111111111111101100","000000000000001001","111111111111101111","000000000000000001","000000000000000011","000000000000010010","000000000000010001","111111111111110011","000000000000000000","111111111111111100","000000000000000001","000000000000001101","000000000000001001","111111111111110101","111111111111110011","000000000000000010","000000000000000100","000000000000000100","111111111111111100","111111111111110100","111111111111111110","111111111111110011","111111111111110000","000000000000000100","000000000000000111","000000000000010011","000000000000001001","111111111111110000","111111111111111010","111111111111111101","000000000000001110","111111111111111011","111111111111110111","111111111111101110","000000000000001100","111111111111101111","000000000000000000","111111111111111110","000000000000001110","000000000000000000","000000000000001001","000000000000000100","000000000000001110","000000000000000000","111111111111110000","111111111111111111","000000000000000111","000000000000000101","111111111111110110","000000000000001011","111111111111101101","111111111111110001","111111111111101110","111111111111110001","111111111111110110","000000000000000110","000000000000000110","000000000000010011","111111111111110100","000000000000000110","000000000000001000","111111111111110000","000000000000001010","000000000000000101","000000000000001111","000000000000000010","000000000000010001","111111111111111111","000000000000010001","000000000000001001","111111111111101100","111111111111111001","000000000000001000","111111111111101110","111111111111110010","111111111111101110","000000000000000001","000000000000001111","111111111111110100","000000000000010000","111111111111111011","000000000000000000","111111111111111000","000000000000001111","000000000000001011","111111111111110000","111111111111111101","111111111111111011","111111111111110100","111111111111110100","111111111111101110","111111111111101101","000000000000000111","000000000000001110","111111111111111110","000000000000001000","000000000000000110","000000000000001101","000000000000000111","000000000000000111","000000000000010010","000000000000000000","000000000000001011","111111111111110110","000000000000000000","000000000000010010","111111111111111010","000000000000010001","111111111111110110","111111111111110011","111111111111101101"),
("111111111111101101","111111111111110011","111111111111110001","111111111111101111","000000000000000000","000000000000001011","000000000000000100","111111111111111000","111111111111101111","111111111111110010","111111111111111010","111111111111111100","000000000000001011","000000000000001101","000000000000000001","000000000000000001","111111111111111001","000000000000001011","000000000000001011","111111111111111011","000000000000000111","000000000000001011","000000000000000100","111111111111110011","111111111111110111","111111111111110111","000000000000000100","111111111111111101","000000000000001000","111111111111111010","000000000000000100","111111111111101100","111111111111110100","111111111111111011","000000000000000101","111111111111110111","000000000000001010","111111111111111101","000000000000001000","111111111111110010","000000000000000010","000000000000000111","000000000000001110","000000000000000101","000000000000000011","111111111111110000","111111111111110001","111111111111110100","000000000000000000","111111111111101101","000000000000001110","111111111111110011","111111111111110001","111111111111110010","111111111111101110","111111111111111000","111111111111110011","111111111111101110","111111111111101101","000000000000010011","111111111111111001","000000000000001101","000000000000010011","111111111111111000","111111111111110001","000000000000000001","111111111111101110","000000000000001111","111111111111110000","000000000000000000","000000000000000010","000000000000000111","111111111111111011","000000000000000100","111111111111111001","111111111111111111","000000000000001111","000000000000001011","000000000000000010","000000000000001010","000000000000000011","111111111111111111","000000000000000001","111111111111111100","111111111111110111","111111111111110010","111111111111111011","111111111111111010","000000000000000111","111111111111110111","000000000000001101","111111111111101101","111111111111101101","111111111111101111","000000000000010010","111111111111110010","111111111111111101","000000000000000000","111111111111101101","000000000000001000","111111111111110101","000000000000000110","111111111111111011","111111111111110100","111111111111110010","000000000000001011","111111111111111100","000000000000010011","111111111111111110","111111111111111011","000000000000001100","000000000000000101","000000000000001110","000000000000000011","000000000000000100","000000000000000000","000000000000010011","000000000000001000","111111111111110000","000000000000000001","000000000000000001","111111111111111001","000000000000010001","000000000000010001","000000000000001110","111111111111111011","000000000000000101","000000000000000000"),
("111111111111110101","000000000000001000","000000000000010011","111111111111111011","000000000000010100","000000000000010010","000000000000010000","111111111111101111","000000000000001110","111111111111101101","111111111111110111","000000000000010010","111111111111111110","111111111111111111","111111111111110101","000000000000010001","000000000000001010","111111111111110110","111111111111111010","000000000000000000","111111111111101100","111111111111111101","111111111111111011","111111111111110111","000000000000001000","000000000000001110","111111111111101101","111111111111101111","111111111111110011","111111111111111110","111111111111110011","000000000000000000","111111111111110110","000000000000010001","111111111111110011","000000000000001100","000000000000000111","111111111111101101","111111111111101111","111111111111111100","000000000000001111","000000000000010100","000000000000001000","111111111111110100","000000000000000000","000000000000001100","111111111111101110","000000000000010001","000000000000000011","000000000000000010","000000000000010000","000000000000000110","111111111111111000","000000000000001100","000000000000010000","000000000000001110","111111111111101101","111111111111110101","000000000000010011","000000000000000010","000000000000000010","111111111111111110","000000000000010000","111111111111101111","000000000000001001","000000000000000001","111111111111111000","111111111111101111","000000000000000101","111111111111111011","000000000000000011","111111111111110100","000000000000010011","000000000000010000","111111111111111010","000000000000001101","111111111111111100","000000000000001110","111111111111110111","000000000000000000","111111111111110000","000000000000000100","111111111111111100","111111111111110001","111111111111101100","000000000000001100","000000000000001011","000000000000000000","111111111111111011","111111111111110011","000000000000010000","111111111111111101","111111111111101111","000000000000000110","111111111111110010","000000000000010000","000000000000001001","000000000000001100","111111111111110101","111111111111101100","111111111111111110","111111111111110001","111111111111111001","000000000000010000","111111111111101111","000000000000001001","000000000000000010","000000000000000010","111111111111111010","000000000000001001","000000000000000000","111111111111110010","111111111111111111","111111111111111001","000000000000010001","000000000000001011","111111111111101111","111111111111111001","000000000000001100","111111111111111000","111111111111111111","000000000000001110","000000000000001101","000000000000010001","000000000000000110","000000000000001010","000000000000010000","111111111111110110"),
("000000000000000110","111111111111111111","000000000000000100","111111111111110000","111111111111111000","000000000000000001","000000000000000100","000000000000000001","111111111111111010","000000000000001101","000000000000001111","111111111111110010","111111111111110001","000000000000010011","000000000000010011","111111111111111001","111111111111110100","000000000000000011","000000000000001000","000000000000000000","000000000000000110","111111111111110110","111111111111110001","111111111111101100","111111111111101101","111111111111111110","000000000000001111","000000000000001111","111111111111111100","111111111111110101","111111111111101101","000000000000010100","000000000000000011","111111111111101101","111111111111110001","111111111111111111","000000000000001001","000000000000001111","111111111111111011","111111111111110010","111111111111110111","000000000000001010","111111111111110111","000000000000001110","000000000000001110","000000000000000010","111111111111110000","000000000000000100","111111111111111010","000000000000001010","000000000000001000","000000000000001000","000000000000010000","111111111111110100","111111111111111110","111111111111111110","000000000000000010","111111111111110100","000000000000000101","111111111111101101","000000000000000001","000000000000001111","111111111111110110","000000000000010001","111111111111110010","111111111111111100","000000000000010010","111111111111111000","111111111111110011","111111111111101110","000000000000010001","000000000000000101","111111111111111110","111111111111111110","111111111111111101","111111111111111010","000000000000001001","111111111111111110","111111111111110000","111111111111110010","111111111111111101","111111111111111100","111111111111111011","111111111111110000","111111111111111111","111111111111110010","000000000000000011","111111111111111011","111111111111110011","111111111111111111","111111111111110000","111111111111111110","111111111111111011","000000000000000100","000000000000001001","111111111111110000","111111111111111100","000000000000000000","000000000000001101","000000000000001010","000000000000010010","000000000000000111","000000000000000000","111111111111111101","000000000000001010","000000000000000000","000000000000000000","111111111111111000","111111111111111000","000000000000010010","000000000000001001","111111111111110111","000000000000000110","000000000000010011","000000000000010011","000000000000010010","111111111111111011","111111111111110101","000000000000000000","111111111111110001","000000000000001011","000000000000000101","111111111111110111","111111111111111101","000000000000000010","000000000000000101","111111111111111000","111111111111110001"),
("000000000000001101","000000000000000110","111111111111110111","111111111111110101","000000000000001000","000000000000000001","000000000000000101","111111111111110111","000000000000000000","000000000000001110","111111111111101100","111111111111110001","000000000000001101","000000000000000110","000000000000000100","111111111111111110","000000000000001111","000000000000000000","000000000000001011","111111111111110111","111111111111101101","000000000000010000","000000000000000000","111111111111110111","111111111111110000","000000000000010001","000000000000001100","111111111111111110","000000000000010000","111111111111111100","111111111111111110","000000000000001001","111111111111111100","000000000000000011","111111111111110000","111111111111110000","111111111111110110","000000000000001011","000000000000001101","000000000000001000","111111111111110001","000000000000010001","111111111111111110","111111111111111100","111111111111110011","000000000000001000","000000000000000011","000000000000010001","111111111111110111","111111111111111100","000000000000001001","111111111111110111","111111111111110111","000000000000001000","000000000000001100","000000000000000001","000000000000000000","000000000000010011","000000000000001111","000000000000010001","000000000000010000","111111111111111001","000000000000010000","000000000000000011","111111111111101100","111111111111110001","000000000000000101","000000000000001010","111111111111110110","111111111111110100","000000000000001010","000000000000001010","111111111111111011","111111111111111010","111111111111110100","000000000000001101","111111111111110001","000000000000001101","111111111111111011","000000000000010011","000000000000000010","111111111111110011","000000000000001000","000000000000001011","000000000000010010","111111111111111011","111111111111101100","111111111111110110","000000000000001111","111111111111111101","111111111111111111","111111111111110110","000000000000000011","000000000000001011","111111111111101100","000000000000010010","111111111111110000","111111111111101110","000000000000001010","000000000000010001","000000000000001000","111111111111101110","000000000000010011","111111111111111000","000000000000001110","000000000000000111","000000000000001110","111111111111111110","000000000000010100","000000000000000101","000000000000001110","000000000000000000","111111111111111011","111111111111111110","000000000000001011","000000000000010011","000000000000001001","111111111111110001","111111111111101111","111111111111111100","111111111111111011","000000000000001001","000000000000000011","111111111111110011","000000000000001010","000000000000000000","111111111111101110","000000000000000100"),
("111111111111110011","000000000000000111","111111111111110010","111111111111111001","111111111111111101","000000000000000001","000000000000000110","111111111111111111","111111111111101101","111111111111101100","111111111111111101","111111111111101110","000000000000010100","000000000000000010","000000000000001010","000000000000010010","000000000000001001","000000000000010011","000000000000000000","000000000000010001","111111111111110101","111111111111111111","000000000000001000","111111111111110101","000000000000000010","111111111111111111","000000000000001010","111111111111110000","111111111111110011","000000000000001110","000000000000010000","000000000000001001","000000000000000011","000000000000001010","111111111111111001","111111111111110001","111111111111111111","111111111111110111","000000000000001101","000000000000000101","000000000000001110","000000000000000101","111111111111110000","111111111111111001","111111111111110011","111111111111111010","000000000000001111","111111111111110101","111111111111111101","111111111111110110","111111111111110001","000000000000000101","111111111111110111","111111111111111110","000000000000000000","000000000000001101","000000000000010001","111111111111101100","000000000000000111","000000000000001101","111111111111101101","000000000000010000","111111111111110111","111111111111101100","111111111111111010","000000000000000100","111111111111101111","000000000000000011","000000000000010000","000000000000000000","000000000000000010","111111111111101110","111111111111111010","000000000000000001","111111111111101110","111111111111110011","111111111111110010","000000000000000111","111111111111110010","111111111111111010","000000000000000011","111111111111111001","111111111111110100","111111111111110110","000000000000010011","111111111111101111","111111111111110000","000000000000001100","111111111111110001","111111111111111011","000000000000000100","111111111111110100","000000000000000100","000000000000001100","111111111111111011","111111111111110111","000000000000000111","111111111111110001","111111111111111110","111111111111111011","111111111111101101","111111111111110101","111111111111110110","111111111111110111","111111111111111001","000000000000000111","000000000000000000","000000000000000001","111111111111101111","000000000000000001","111111111111111111","111111111111111100","000000000000010100","111111111111111011","000000000000001000","000000000000001010","111111111111111101","111111111111111101","111111111111101111","111111111111111000","111111111111110111","111111111111110011","111111111111110100","000000000000000000","111111111111110010","000000000000000110","000000000000000100","111111111111101111"),
("111111111111111111","111111111111111111","111111111111111101","000000000000001001","000000000000000000","000000000000000110","111111111111110001","000000000000000000","000000000000000001","111111111111101111","111111111111110101","000000000000001011","000000000000000011","000000000000001010","000000000000000011","111111111111101101","000000000000001011","000000000000001001","111111111111101110","000000000000001010","111111111111111110","111111111111110100","000000000000010001","111111111111101110","000000000000000101","000000000000001010","000000000000000110","111111111111111000","111111111111111101","111111111111111011","111111111111110110","000000000000001010","111111111111110110","111111111111101101","111111111111101100","000000000000000111","111111111111111010","111111111111111000","000000000000000000","111111111111110011","111111111111110010","000000000000010000","000000000000000100","000000000000000111","000000000000001100","111111111111111011","111111111111110010","000000000000010011","111111111111110100","000000000000000101","111111111111110001","000000000000000001","000000000000000011","111111111111111000","000000000000010000","111111111111110000","111111111111110101","000000000000001101","000000000000001111","111111111111110111","000000000000000111","000000000000001110","000000000000010001","000000000000000000","111111111111110001","000000000000001000","111111111111110111","111111111111111001","111111111111110000","111111111111110110","000000000000000100","111111111111111101","111111111111110101","111111111111111010","111111111111111000","111111111111111110","111111111111101110","111111111111110011","000000000000001011","000000000000001101","111111111111110010","111111111111110101","000000000000000111","000000000000001001","000000000000000100","111111111111110111","000000000000000011","111111111111110100","111111111111111101","111111111111110000","000000000000001111","000000000000000010","111111111111110101","111111111111110110","000000000000000111","000000000000001101","111111111111111011","111111111111111011","000000000000000101","000000000000001110","000000000000000101","111111111111110001","111111111111110110","000000000000010001","111111111111110010","000000000000001110","000000000000000100","000000000000000100","000000000000010001","111111111111101101","000000000000000000","000000000000001010","000000000000000010","000000000000000000","000000000000000101","111111111111111111","111111111111101110","111111111111110001","111111111111101110","111111111111111000","000000000000001110","000000000000000000","000000000000000101","000000000000000011","111111111111111000","111111111111111100","000000000000000111","000000000000000101"),
("111111111111111000","111111111111110000","000000000000000100","000000000000001010","111111111111110011","111111111111101110","000000000000010011","111111111111110010","000000000000010001","111111111111110101","111111111111110111","000000000000000010","111111111111111101","111111111111111100","111111111111111011","000000000000001010","111111111111111100","111111111111110111","000000000000001101","000000000000010001","000000000000010001","111111111111110010","111111111111111100","000000000000000010","000000000000000000","111111111111110101","000000000000000101","111111111111111100","111111111111110110","111111111111111010","000000000000010000","111111111111110111","000000000000000100","000000000000000110","111111111111111000","000000000000001101","111111111111110001","111111111111111100","000000000000010100","000000000000001111","111111111111110001","000000000000001011","111111111111110100","111111111111110000","000000000000000001","000000000000000110","000000000000001000","000000000000000100","111111111111110111","111111111111111110","111111111111111000","111111111111111001","000000000000000101","000000000000001011","000000000000001011","000000000000000011","111111111111101101","000000000000000000","000000000000001000","111111111111110100","000000000000010000","111111111111110001","111111111111101100","111111111111111011","000000000000001110","000000000000001010","000000000000000100","000000000000010100","000000000000000111","111111111111111110","111111111111111110","000000000000010000","000000000000010010","111111111111111000","000000000000001100","111111111111110001","111111111111101101","000000000000001100","000000000000001001","000000000000001000","000000000000001100","000000000000010000","111111111111110101","111111111111110101","111111111111110101","111111111111111100","000000000000001010","111111111111111110","111111111111101110","111111111111111100","111111111111111011","111111111111111001","111111111111101101","000000000000000000","000000000000001001","000000000000001011","111111111111111110","111111111111101111","111111111111111110","000000000000000000","000000000000010100","111111111111110111","000000000000010011","111111111111110110","111111111111101100","111111111111110101","111111111111111100","111111111111110100","111111111111110101","111111111111110100","111111111111101111","000000000000010100","000000000000000001","111111111111110011","000000000000000111","111111111111111001","000000000000001101","111111111111111111","000000000000000101","000000000000000110","111111111111101101","111111111111111011","000000000000000110","000000000000010000","000000000000001000","111111111111110010","000000000000000011","000000000000000000"),
("111111111111110010","111111111111111011","000000000000001011","000000000000010100","000000000000001010","000000000000001000","111111111111110010","111111111111101110","000000000000001001","000000000000001100","111111111111110001","000000000000001101","000000000000001011","000000000000000011","000000000000000000","000000000000010011","111111111111101100","111111111111101111","000000000000000111","000000000000000001","111111111111101100","000000000000001100","000000000000000100","111111111111111010","000000000000001000","111111111111101101","000000000000000001","111111111111111111","000000000000000011","000000000000010010","000000000000001110","000000000000000010","111111111111101101","000000000000000010","111111111111111100","111111111111111011","000000000000000010","000000000000000001","000000000000010100","000000000000001111","000000000000000100","111111111111111011","111111111111101111","000000000000001010","111111111111101101","000000000000001001","111111111111110000","111111111111111000","111111111111110100","111111111111110101","000000000000010011","000000000000010100","111111111111101110","000000000000000001","000000000000001011","000000000000001100","000000000000001110","111111111111111100","000000000000010001","111111111111111110","111111111111111000","111111111111110011","111111111111111100","111111111111110110","111111111111110001","111111111111110001","111111111111110111","111111111111110010","000000000000000001","111111111111110111","000000000000010000","111111111111111100","000000000000001110","111111111111101100","000000000000000000","000000000000001111","111111111111101110","111111111111110000","000000000000001110","000000000000000000","000000000000001001","111111111111111100","111111111111110000","111111111111101100","000000000000000110","111111111111110101","111111111111110001","111111111111111010","000000000000001111","111111111111110101","000000000000000000","000000000000001011","111111111111101101","111111111111110101","111111111111101110","111111111111111001","000000000000000010","000000000000000110","000000000000010001","111111111111111000","000000000000000000","111111111111111011","000000000000010010","000000000000001010","000000000000000100","111111111111110001","111111111111110110","000000000000001000","000000000000001000","000000000000010100","111111111111111110","000000000000001101","111111111111110000","111111111111101101","000000000000001111","000000000000001010","111111111111110100","111111111111111000","000000000000001110","000000000000001110","111111111111110100","111111111111111101","111111111111111111","000000000000000100","111111111111111100","000000000000001011","111111111111110010","111111111111111001"),
("000000000000001110","111111111111111111","111111111111111000","000000000000010000","111111111111111110","000000000000000001","000000000000001111","000000000000000110","000000000000000000","000000000000001101","000000000000001011","000000000000000001","000000000000000000","111111111111101111","000000000000000110","000000000000001101","000000000000010001","000000000000010000","000000000000001011","000000000000001110","000000000000001010","111111111111101100","111111111111111110","000000000000001001","111111111111101111","000000000000000100","111111111111111100","111111111111111110","111111111111111100","111111111111110111","111111111111111100","111111111111110011","000000000000000000","000000000000010000","111111111111110010","000000000000001111","000000000000010100","000000000000001000","111111111111111010","111111111111111110","000000000000010001","000000000000010000","000000000000000010","000000000000000001","000000000000000001","000000000000010000","111111111111111000","111111111111101110","000000000000000011","000000000000010001","000000000000001111","111111111111110111","000000000000001100","000000000000010011","111111111111110111","111111111111110111","111111111111111001","000000000000000101","111111111111110110","111111111111101110","111111111111110000","000000000000000110","111111111111110000","111111111111111001","000000000000010100","000000000000001100","111111111111101110","000000000000010011","111111111111101100","000000000000000000","000000000000000001","000000000000000101","111111111111110001","111111111111101110","000000000000001000","111111111111110001","111111111111110100","111111111111110000","111111111111101100","000000000000000101","000000000000001011","111111111111101111","000000000000000111","000000000000000011","000000000000000110","111111111111110010","000000000000010001","000000000000000111","111111111111111110","000000000000001001","111111111111111010","111111111111101111","000000000000000101","111111111111101111","000000000000000100","000000000000001100","111111111111101100","000000000000001000","000000000000001010","000000000000001000","000000000000010001","000000000000010010","111111111111111101","111111111111101101","000000000000001010","111111111111110101","111111111111111100","000000000000001010","000000000000000010","111111111111111010","111111111111111000","000000000000001110","111111111111101101","000000000000000011","000000000000001110","000000000000000110","111111111111111011","000000000000000100","111111111111111001","000000000000010011","000000000000010011","111111111111111100","000000000000000100","000000000000000110","111111111111110010","111111111111110100","111111111111110000","111111111111111111"),
("111111111111110000","000000000000000000","000000000000000000","000000000000001111","111111111111111111","000000000000000110","000000000000000001","111111111111110101","111111111111111011","000000000000010100","111111111111110111","000000000000001100","000000000000010000","111111111111110110","111111111111111101","111111111111101101","111111111111110110","000000000000000010","000000000000001101","000000000000000000","000000000000001100","111111111111110111","000000000000001001","000000000000000110","000000000000001010","000000000000000010","000000000000010011","111111111111111111","111111111111110110","000000000000010100","000000000000001100","111111111111110001","111111111111110011","111111111111110001","000000000000010010","111111111111110101","111111111111110100","000000000000000000","000000000000000101","000000000000010011","111111111111111111","111111111111111010","111111111111101110","000000000000001110","111111111111111101","111111111111111100","000000000000010000","111111111111110110","000000000000001110","111111111111111011","000000000000001100","111111111111111000","000000000000000101","111111111111111011","111111111111101111","000000000000001110","000000000000000100","111111111111110100","000000000000010000","000000000000001000","111111111111110111","000000000000001011","000000000000001110","000000000000010100","111111111111111010","000000000000010010","000000000000001101","000000000000000100","000000000000001100","000000000000001010","000000000000001110","000000000000000000","000000000000010010","111111111111111011","000000000000001101","111111111111110110","000000000000001010","000000000000000000","111111111111110010","111111111111101110","000000000000001111","111111111111111010","000000000000000001","000000000000000111","111111111111101111","000000000000000000","000000000000010001","111111111111111110","111111111111110100","111111111111101110","000000000000000001","000000000000001110","000000000000010100","000000000000000011","111111111111111000","111111111111111111","111111111111111101","000000000000000010","111111111111110000","111111111111111001","111111111111110010","000000000000000100","000000000000001000","111111111111111011","111111111111110110","111111111111111100","111111111111110001","000000000000001111","111111111111110111","000000000000001011","111111111111111101","111111111111110101","111111111111101100","000000000000000011","111111111111110110","111111111111110011","000000000000000000","111111111111111100","111111111111101100","111111111111111010","111111111111101111","111111111111110011","000000000000010001","111111111111111001","000000000000001000","111111111111111101","111111111111101111","111111111111110111"),
("111111111111110010","000000000000001000","111111111111101110","111111111111110100","111111111111110000","111111111111110010","111111111111101110","000000000000001000","111111111111101100","111111111111111001","111111111111110100","000000000000000110","111111111111101111","000000000000010001","111111111111101111","111111111111110011","000000000000001001","111111111111111010","000000000000001010","000000000000001011","000000000000000100","111111111111101111","000000000000000101","111111111111110101","111111111111111011","111111111111110010","111111111111111001","000000000000010100","000000000000001001","000000000000000000","000000000000010001","000000000000000010","111111111111111111","000000000000010001","111111111111110000","000000000000001011","111111111111111011","000000000000000010","000000000000000110","111111111111110101","111111111111111100","000000000000001010","000000000000001011","000000000000000010","111111111111111101","111111111111111000","111111111111111001","111111111111110100","000000000000000000","111111111111111101","000000000000000000","000000000000001110","111111111111110000","000000000000001000","111111111111111010","111111111111111011","000000000000000100","111111111111101110","111111111111111010","111111111111111110","111111111111111101","111111111111110110","000000000000001011","000000000000000011","111111111111110100","000000000000010000","111111111111110000","000000000000001100","000000000000010000","000000000000000000","000000000000001011","000000000000000000","000000000000010011","111111111111110110","111111111111111111","111111111111110100","000000000000000011","000000000000000000","000000000000010010","000000000000000011","111111111111110100","111111111111110101","000000000000010011","000000000000000101","000000000000001111","000000000000001110","000000000000001110","000000000000001011","000000000000010011","000000000000001000","000000000000001001","111111111111111100","000000000000000000","000000000000000111","000000000000001000","000000000000001110","000000000000000001","000000000000001101","000000000000001011","000000000000001101","000000000000000000","000000000000001111","000000000000000100","000000000000000011","000000000000000110","000000000000001001","111111111111111000","000000000000001100","111111111111110100","000000000000000010","111111111111101100","000000000000001001","111111111111101101","000000000000010001","000000000000000010","000000000000000000","000000000000001000","000000000000000001","000000000000001101","111111111111111001","111111111111101110","111111111111101101","111111111111111100","000000000000001010","000000000000000000","000000000000000000","111111111111110011","111111111111111001"),
("000000000000000111","000000000000010010","000000000000001000","111111111111110011","000000000000001100","000000000000010000","000000000000001001","111111111111111100","000000000000000110","000000000000001111","111111111111111000","000000000000011101","111111111111111110","000000000000001101","000000000000000110","000000000000000001","000000000000001011","111111111111111101","111111111111101111","111111111111110001","111111111111110000","111111111111101110","000000000000000101","111111111111111111","000000000000000111","000000000000000001","000000000000001000","000000000000001000","111111111111111100","000000000000000001","111111111111101111","000000000000010110","000000000000000000","000000000000100010","000000000000000000","111111111111111000","000000000000001111","000000000000000001","000000000000000010","111111111111111001","000000000000001110","000000000000100001","111111111111111010","000000000000001000","111111111111101000","000000000000000101","000000000000000000","111111111111111101","111111111111101101","000000000000001110","111111111111111010","000000000000000101","000000000000011001","111111111111110101","000000000000000110","111111111111101101","000000000000000000","000000000000000001","111111111111110001","000000000000000110","111111111111110100","000000000000001000","111111111111111010","000000000000001100","000000000000000001","000000000000011010","111111111111110101","000000000000001101","111111111111111100","111111111111111011","111111111111110100","000000000000010110","111111111111110000","000000000000000001","000000000000000110","111111111111110101","000000000000000010","000000000000000001","111111111111111100","111111111111101110","111111111111110010","111111111111110111","111111111111011110","000000000000010000","111111111111101000","000000000000010100","111111111111101110","000000000000011011","111111111111111011","000000000000001010","111111111111111110","000000000000000001","000000000000010011","000000000000010100","000000000000000101","000000000000010000","111111111111111111","000000000000000001","000000000000000110","111111111111111111","000000000000010100","000000000000001110","111111111111111100","111111111111101001","111111111111110101","111111111111111000","000000000000001100","000000000000010111","111111111111110111","111111111111101000","000000000000000010","000000000000000100","111111111111111111","000000000000000100","000000000000001101","000000000000010110","000000000000010010","111111111111111011","111111111111111000","111111111111101110","111111111111111001","000000000000000110","000000000000011000","000000000000001011","111111111111110010","111111111111111011","111111111111111000","111111111111110010"),
("000000000000001110","000000000000001110","111111111111101011","111111111111111001","000000000000000000","000000000000001010","000000000000001111","111111111111101100","000000000000000000","000000000000000110","000000000000001000","000000000000010010","000000000000001010","111111111111111010","000000000000001100","111111111111111101","111111111111110000","111111111111110101","111111111111111111","000000000000000110","000000000000010001","111111111111111111","111111111111110011","111111111111101110","000000000000001011","000000000000000000","000000000000000000","000000000000011010","111111111111111100","000000000000000000","000000000000000001","000000000000000001","000000000000000111","111111111111111110","111111111111110111","000000000000001100","000000000000001101","111111111111110000","111111111111101110","111111111111110010","000000000000001000","000000000000010010","111111111111111000","000000000000000011","111111111111110011","000000000000010001","111111111111111101","000000000000001101","000000000000001010","000000000000010101","111111111111111000","000000000000001000","111111111111110111","111111111111100010","000000000000000100","000000000000001010","000000000000000000","000000000000000111","000000000000000100","000000000000000000","000000000000010100","000000000000000011","000000000000000000","111111111111101111","111111111111111100","000000000000000000","000000000000010000","111111111111111100","111111111111100101","000000000000001001","000000000000010110","000000000000000000","000000000000000010","111111111111110001","000000000000000110","000000000000001001","111111111111101011","000000000000011001","111111111111101100","111111111111111110","111111111111111001","111111111111100101","111111111111111000","111111111111111111","111111111111110110","111111111111101111","000000000000000010","000000000000001111","000000000000011110","111111111111111011","000000000000011110","111111111111111101","000000000000001010","111111111111111101","111111111111110111","111111111111110100","111111111111111110","111111111111111100","111111111111111001","000000000000001111","111111111111111101","000000000000100000","000000000000000011","111111111111101011","111111111111110100","111111111111110001","111111111111110011","000000000000010001","111111111111111100","111111111111101010","111111111111111001","111111111111111111","000000000000001001","000000000000000101","000000000000000100","000000000000010010","000000000000010110","111111111111111100","000000000000010001","111111111111111110","000000000000001110","000000000000000101","000000000000010000","111111111111101101","000000000000000111","000000000000001000","000000000000001000","111111111111110111"),
("111111111111110111","111111111111011101","111111111111111110","000000000000000111","000000000000000011","000000000000001110","000000000000011010","111111111111111010","000000000000001100","111111111111110000","000000000000001101","111111111111111011","111111111111110111","111111111111111010","000000000000001100","000000000000000000","111111111111110111","000000000000000100","000000000000000011","000000000000000000","111111111111111000","000000000000000101","111111111111110000","000000000000000000","111111111111111001","000000000000001111","000000000000010001","000000000000000010","111111111111101101","111111111111110001","111111111111111010","000000000000000101","111111111111111011","000000000000001110","000000000000001010","111111111111110000","000000000000010101","111111111111110010","111111111111110100","000000000000001011","111111111111110000","111111111111101101","000000000000010011","000000000000010111","111111111111111010","111111111111101110","111111111111111110","000000000000010011","111111111111110011","111111111111101011","000000000000000100","111111111111111000","000000000000001110","000000000000001111","000000000000010011","000000000000000111","111111111111101100","000000000000000011","111111111111101010","000000000000010100","111111111111111001","000000000000000000","000000000000000111","000000000000000100","000000000000000111","111111111111101100","111111111111110110","111111111111110111","000000000000000110","111111111111110100","000000000000010110","000000000000010101","000000000000000100","000000000000001001","000000000000000010","111111111111111101","000000000000000100","000000000000001111","111111111111101010","111111111111111011","000000000000000111","111111111111111011","000000000000000101","000000000000000101","000000000000001110","111111111111111100","000000000000010011","000000000000000110","000000000000001011","000000000000010011","000000000000001000","111111111111110110","111111111111111011","000000000000011011","111111111111111000","000000000000000110","000000000000000110","000000000000011011","111111111111100110","000000000000000001","000000000000000011","000000000000001011","000000000000000110","111111111111111011","000000000000010100","000000000000001110","000000000000000000","000000000000001001","000000000000001110","111111111111110001","111111111111110011","111111111111111100","111111111111110011","000000000000000110","000000000000010001","000000000000011111","000000000000010000","000000000000010100","111111111111110100","111111111111111100","000000000000010100","111111111111110001","000000000000010111","000000000000001011","000000000000000000","111111111111101001","111111111111110110","111111111111110011"),
("111111111111110100","000000000000000110","111111111111101110","000000000000010010","111111111111101001","000000000000001000","000000000000010010","111111111111110011","111111111111110011","000000000000001101","111111111111111110","000000000000001011","111111111111110111","111111111111110011","111111111111101100","111111111111110110","000000000000000010","000000000000000011","111111111111110010","111111111111110010","000000000000000100","000000000000000000","111111111111101000","111111111111111111","000000000000000110","000000000000001101","000000000000010010","000000000000010100","000000000000010011","111111111111111110","000000000000000000","111111111111101110","111111111111111101","111111111111110100","000000000000000000","111111111111111011","000000000000001101","000000000000001101","000000000000001000","000000000000001101","000000000000001000","000000000000010000","000000000000001010","000000000000010100","000000000000001101","111111111111111111","000000000000000001","000000000000010001","000000000000000000","000000000000001110","000000000000001001","111111111111111001","111111111111111110","000000000000000010","000000000000000011","111111111111111001","000000000000001000","000000000000000111","111111111111111010","000000000000000100","111111111111111000","111111111111110100","000000000000001111","111111111111101110","000000000000001100","111111111111110001","000000000000001111","000000000000001001","000000000000001111","111111111111101101","000000000000000010","111111111111101111","111111111111111001","111111111111101110","111111111111101101","000000000000001111","000000000000010010","000000000000000111","000000000000000000","000000000000010000","111111111111110000","000000000000000010","111111111111110001","111111111111101001","000000000000000110","000000000000000001","000000000000001010","000000000000000001","111111111111111010","111111111111101110","111111111111110110","111111111111111111","111111111111101101","111111111111111110","000000000000001110","111111111111111011","111111111111110111","000000000000001110","111111111111101100","000000000000010011","000000000000001011","111111111111111001","000000000000000000","000000000000000001","111111111111110011","111111111111110000","111111111111111110","000000000000001011","000000000000001100","111111111111110100","111111111111111010","000000000000000101","000000000000000111","111111111111110011","000000000000000100","000000000000001110","000000000000000100","000000000000010010","000000000000000000","000000000000000010","111111111111110111","000000000000001000","111111111111111000","111111111111110101","111111111111111110","111111111111111010","000000000000000110","000000000000001001"),
("111111111111110110","000000000000000101","111111111111110110","000000000000001110","000000000000010010","000000000000000001","111111111111111010","111111111111111010","000000000000000100","000000000000001111","111111111111110001","111111111111101100","000000000000000000","111111111111110011","000000000000001100","000000000000001010","000000000000000110","000000000000001101","111111111111110001","111111111111111000","000000000000001001","000000000000000100","111111111111101110","000000000000001111","111111111111111111","111111111111111111","000000000000000101","111111111111111110","000000000000010100","111111111111111011","000000000000000101","000000000000001000","111111111111110010","111111111111111011","111111111111111111","111111111111110110","000000000000000010","000000000000000101","000000000000001100","111111111111110110","111111111111110100","000000000000001011","111111111111101110","111111111111111110","111111111111111010","000000000000000001","000000000000010011","000000000000001000","000000000000000101","000000000000000101","111111111111111010","111111111111111111","000000000000010000","000000000000010100","111111111111111010","000000000000010011","000000000000000011","000000000000000111","000000000000000011","000000000000001010","111111111111110111","000000000000000110","111111111111111110","111111111111101101","111111111111110111","000000000000001011","000000000000001101","111111111111101111","000000000000000001","111111111111111101","000000000000001010","111111111111111011","000000000000000000","000000000000001110","000000000000001001","111111111111111101","111111111111111011","000000000000000010","111111111111110010","111111111111101111","111111111111110011","000000000000000010","000000000000000110","111111111111101111","000000000000010010","111111111111110101","111111111111110110","000000000000001001","000000000000000000","000000000000010000","000000000000010000","111111111111110100","000000000000000101","000000000000001110","111111111111110111","000000000000001010","000000000000010000","000000000000001111","000000000000001000","000000000000000100","111111111111111011","000000000000000111","111111111111110101","111111111111111100","000000000000010010","000000000000010010","000000000000000000","000000000000000011","000000000000000110","000000000000000000","111111111111101110","111111111111110101","111111111111101101","000000000000010010","111111111111110101","111111111111111100","111111111111101101","111111111111101101","111111111111111010","111111111111111101","000000000000000011","000000000000000111","000000000000000001","000000000000010000","111111111111110010","000000000000010011","000000000000001010","000000000000001010"),
("000000000000000101","000000000000001010","000000000000000001","000000000000001111","111111111111111110","111111111111111111","111111111111111010","111111111111101100","000000000000000011","111111111111111110","111111111111110110","000000000000000000","000000000000000100","111111111111110001","111111111111111100","000000000000001111","111111111111111000","111111111111101111","000000000000000011","000000000000010010","111111111111111010","111111111111111000","111111111111111001","111111111111110010","111111111111111011","000000000000000010","000000000000000000","111111111111110011","111111111111111101","000000000000001010","111111111111111010","000000000000001101","111111111111110001","000000000000001000","000000000000001101","111111111111111010","000000000000000001","000000000000001000","000000000000010010","111111111111111010","000000000000000000","111111111111110110","111111111111101111","111111111111111111","000000000000000111","000000000000001000","000000000000001101","111111111111111001","000000000000000011","111111111111111000","111111111111101110","000000000000001001","111111111111101110","000000000000010010","111111111111111010","000000000000010001","000000000000000100","111111111111101101","000000000000000100","000000000000000100","000000000000001110","111111111111111101","000000000000000100","111111111111101111","000000000000000000","000000000000000000","000000000000000100","000000000000000100","111111111111110001","000000000000000110","111111111111110001","111111111111111101","000000000000000010","111111111111111000","111111111111111110","111111111111110000","000000000000010000","000000000000000111","111111111111111001","000000000000000011","111111111111110000","000000000000001110","000000000000001011","111111111111110010","000000000000000011","000000000000010100","000000000000001101","000000000000000111","000000000000000111","000000000000000100","111111111111101101","111111111111111000","000000000000000100","000000000000001010","111111111111110000","000000000000000110","111111111111101100","111111111111101100","000000000000010000","111111111111111100","111111111111110001","000000000000001100","111111111111101100","000000000000000101","111111111111101110","000000000000001111","000000000000000000","000000000000000101","111111111111111110","000000000000001110","000000000000001100","111111111111101101","000000000000000011","000000000000010100","000000000000010010","111111111111111100","000000000000000000","111111111111101111","000000000000000111","000000000000000100","111111111111111011","111111111111101101","111111111111110100","111111111111101111","000000000000000000","111111111111110000","000000000000000011","111111111111110001"),
("000000000000000111","111111111111101101","111111111111111111","000000000000000000","000000000000000111","000000000000000100","000000000000001010","000000000000001110","111111111111110111","000000000000000000","111111111111111110","000000000000010000","000000000000001010","000000000000001010","111111111111111110","000000000000001110","111111111111110001","000000000000000101","000000000000000110","000000000000001101","111111111111110011","111111111111111110","111111111111110011","000000000000001000","000000000000001001","000000000000001111","000000000000010000","000000000000000011","111111111111110110","000000000000000000","111111111111101100","111111111111111010","000000000000001100","000000000000000010","000000000000010011","111111111111111001","111111111111110001","111111111111111000","000000000000010010","000000000000001001","000000000000001111","111111111111111101","111111111111110011","111111111111111001","000000000000001001","000000000000000010","000000000000000111","000000000000001000","111111111111110001","000000000000001001","111111111111111111","000000000000010000","111111111111110101","000000000000010100","000000000000010100","111111111111111011","111111111111111101","000000000000000101","111111111111110111","000000000000001000","111111111111101100","000000000000001100","000000000000000110","111111111111111010","111111111111111000","111111111111101110","000000000000000101","111111111111111000","111111111111111011","000000000000001011","111111111111111100","000000000000001000","000000000000000010","111111111111111001","111111111111111000","111111111111101110","000000000000000000","111111111111111000","111111111111110010","111111111111110110","111111111111111010","000000000000001100","111111111111110101","000000000000000010","111111111111101101","000000000000000101","000000000000000110","111111111111101101","111111111111111010","111111111111110001","111111111111111001","111111111111110111","000000000000000111","111111111111110011","000000000000010001","000000000000001000","000000000000010011","111111111111111001","111111111111110011","000000000000001101","000000000000001010","111111111111111111","111111111111110011","111111111111110101","111111111111110001","111111111111110110","000000000000001101","000000000000000010","111111111111111111","111111111111110001","000000000000001010","000000000000001010","111111111111111110","111111111111110110","111111111111111011","000000000000000010","000000000000000000","000000000000000001","111111111111101100","111111111111101101","000000000000000001","000000000000000101","111111111111110101","000000000000001100","111111111111110100","000000000000000100","000000000000001010","000000000000010010"),
("111111111111111010","000000000000000001","000000000000000010","000000000000000000","000000000000000100","000000000000000101","000000000000000100","000000000000000001","000000000000000101","111111111111110011","000000000000000011","000000000000000010","111111111111110000","000000000000000100","000000000000001101","000000000000010100","000000000000001100","111111111111101101","000000000000010010","111111111111101101","111111111111110101","111111111111110110","111111111111101110","111111111111101100","000000000000001010","000000000000000011","111111111111111100","111111111111110111","000000000000001001","111111111111110100","111111111111111011","111111111111101101","000000000000000111","000000000000000000","111111111111110100","000000000000001110","000000000000000011","000000000000010011","000000000000000000","000000000000000111","111111111111111010","111111111111110111","111111111111110110","111111111111101110","000000000000001000","000000000000000100","000000000000001010","000000000000001010","000000000000001011","000000000000000101","000000000000001111","000000000000010001","111111111111110100","111111111111111111","000000000000001011","111111111111110110","111111111111111001","111111111111110111","000000000000010000","111111111111110101","111111111111110100","111111111111101110","000000000000000000","000000000000010010","111111111111111010","000000000000000011","000000000000000011","111111111111101101","111111111111111110","111111111111111100","000000000000001111","111111111111110110","000000000000001101","000000000000001101","000000000000001111","000000000000000010","000000000000000010","111111111111110101","111111111111110101","000000000000001011","000000000000001000","111111111111111101","111111111111111101","000000000000001101","111111111111110110","111111111111110100","111111111111111011","000000000000010010","000000000000000110","000000000000001010","111111111111110111","111111111111101101","000000000000010010","111111111111110000","111111111111111111","000000000000000000","000000000000010000","000000000000010011","000000000000000110","000000000000010100","000000000000001100","000000000000001010","111111111111110100","000000000000000110","111111111111111110","000000000000000101","111111111111110111","000000000000010001","000000000000000011","111111111111111011","000000000000000000","111111111111110111","111111111111111011","000000000000000000","000000000000001101","000000000000001011","111111111111111000","000000000000001000","000000000000001100","000000000000001011","111111111111110110","000000000000001000","000000000000010001","000000000000010100","111111111111110010","000000000000000000","111111111111111000","111111111111111011"),
("111111111111110011","111111111111110111","000000000000000110","111111111111110110","111111111111111101","111111111111110100","111111111111111100","111111111111110110","111111111111101101","111111111111101111","000000000000001000","000000000000010100","000000000000000001","000000000000001110","000000000000001010","000000000000000100","111111111111111001","111111111111110101","000000000000000010","000000000000010001","000000000000010100","111111111111111101","111111111111111101","000000000000001101","111111111111111111","111111111111111000","000000000000010100","111111111111111111","111111111111110111","000000000000000010","000000000000001000","000000000000000100","000000000000001100","111111111111101101","111111111111110000","000000000000000001","000000000000010010","111111111111111101","111111111111110000","000000000000000001","000000000000001011","111111111111110001","000000000000001110","000000000000000010","111111111111110100","000000000000000110","000000000000001011","111111111111110010","000000000000000010","000000000000000000","111111111111101101","111111111111101110","111111111111111100","000000000000001100","111111111111101110","000000000000001010","000000000000000110","111111111111110110","000000000000001111","000000000000000000","000000000000001010","000000000000000000","111111111111110001","000000000000000011","111111111111110111","000000000000010001","000000000000001111","111111111111110101","111111111111101111","111111111111101111","111111111111110111","000000000000001001","111111111111111011","000000000000000101","000000000000001110","111111111111101110","111111111111110010","111111111111111011","000000000000010000","111111111111110111","111111111111111110","000000000000001010","111111111111111010","111111111111110111","111111111111111010","000000000000010011","000000000000001101","111111111111110010","000000000000000000","111111111111110111","000000000000000111","111111111111111011","111111111111110010","111111111111110100","000000000000010001","000000000000010011","000000000000001011","000000000000000110","111111111111111010","111111111111101101","111111111111110101","000000000000001000","000000000000000001","111111111111110000","000000000000000000","000000000000010001","000000000000000000","000000000000001111","000000000000000101","111111111111110100","111111111111111010","000000000000001101","000000000000001011","111111111111110000","111111111111111010","000000000000010011","000000000000001001","111111111111111110","000000000000000101","000000000000001001","111111111111110111","000000000000001001","000000000000000001","000000000000001011","111111111111110010","000000000000001011","111111111111110001","000000000000001001"),
("111111111111111111","111111111111111011","111111111111111110","000000000000000100","111111111111111101","000000000000000111","111111111111111101","111111111111101110","000000000000001010","111111111111110010","000000000000000001","000000000000001001","000000000000001100","111111111111110010","000000000000010100","111111111111111100","000000000000001110","000000000000001101","111111111111110011","000000000000010001","111111111111111110","111111111111110111","111111111111111000","000000000000000001","111111111111101101","111111111111110011","111111111111101111","111111111111101101","111111111111111101","000000000000010001","111111111111111010","000000000000000111","000000000000001110","000000000000000101","111111111111110101","000000000000001100","000000000000000000","111111111111111000","000000000000010000","000000000000000000","000000000000001011","111111111111110100","000000000000001100","000000000000000000","000000000000001001","111111111111110000","111111111111110011","000000000000000101","000000000000010001","000000000000001000","111111111111101110","000000000000001000","111111111111101110","111111111111110111","000000000000010100","111111111111111111","111111111111110100","000000000000010010","111111111111110011","111111111111111001","000000000000000000","111111111111110000","111111111111101100","000000000000000100","000000000000000111","000000000000000110","000000000000000101","000000000000000110","000000000000001111","000000000000001010","111111111111110110","000000000000001010","111111111111101111","111111111111111111","111111111111101101","111111111111111001","000000000000010100","000000000000010000","000000000000000101","000000000000010100","111111111111101111","000000000000001101","000000000000000010","111111111111101110","111111111111111010","111111111111111101","111111111111111001","000000000000000100","111111111111110010","111111111111101100","000000000000001011","111111111111111110","111111111111111100","111111111111110101","000000000000010001","111111111111111111","111111111111101111","000000000000010000","000000000000010000","000000000000001101","111111111111111111","111111111111111000","111111111111110110","000000000000010100","111111111111101110","111111111111110110","000000000000001111","111111111111110011","000000000000010010","111111111111111001","000000000000000100","000000000000000001","111111111111111111","111111111111110111","000000000000010001","111111111111111110","000000000000001001","111111111111111100","111111111111110010","111111111111101110","000000000000000000","000000000000001101","000000000000000111","000000000000001100","111111111111101111","000000000000010100","111111111111111110","000000000000000000"),
("111111111111111110","111111111111111001","111111111111111011","000000000000000001","111111111111110010","000000000000010000","111111111111110110","111111111111110110","111111111111111011","111111111111110110","000000000000000011","000000000000000101","111111111111101111","000000000000001100","000000000000001001","111111111111110001","111111111111111000","000000000000000000","000000000000000011","111111111111110001","111111111111110100","111111111111101111","000000000000000010","111111111111111011","000000000000000000","111111111111110100","000000000000001010","111111111111111000","000000000000000100","111111111111111001","000000000000000000","000000000000001001","111111111111111111","000000000000010001","000000000000001010","111111111111110111","000000000000000000","111111111111110110","000000000000000101","000000000000000010","111111111111111101","111111111111110101","111111111111111011","000000000000001011","111111111111111001","000000000000000001","000000000000000101","000000000000000001","111111111111111110","111111111111101101","000000000000010010","111111111111111101","111111111111111000","000000000000010011","000000000000000101","000000000000000011","000000000000000100","111111111111110000","111111111111111011","000000000000001011","111111111111101111","000000000000001000","000000000000000000","000000000000001010","111111111111111110","000000000000001001","111111111111111001","111111111111101101","111111111111101100","000000000000000010","111111111111110001","111111111111111010","000000000000000001","111111111111111111","111111111111111101","000000000000000001","000000000000010000","111111111111101110","000000000000001100","000000000000001000","000000000000000010","111111111111111011","111111111111110100","111111111111101100","000000000000000010","000000000000010100","000000000000001010","000000000000000101","111111111111111110","111111111111111011","000000000000001111","111111111111110011","111111111111110101","111111111111110110","000000000000010010","111111111111110011","111111111111110101","111111111111111000","111111111111110111","000000000000000001","000000000000000011","000000000000000101","111111111111110001","000000000000000110","111111111111110110","000000000000001011","000000000000000110","000000000000001101","111111111111111110","000000000000000010","111111111111111100","000000000000001100","111111111111110101","000000000000001011","000000000000000101","111111111111110000","000000000000001101","000000000000000101","000000000000000000","000000000000001000","000000000000000001","111111111111101101","111111111111101110","000000000000001000","000000000000001110","000000000000001101","000000000000001000","000000000000010100"),
("000000000000000000","000000000000010000","111111111111110010","000000000000001001","000000000000000100","111111111111111101","111111111111110100","000000000000001100","111111111111111100","111111111111111111","111111111111110001","111111111111111111","111111111111110010","111111111111111010","000000000000010000","111111111111111001","000000000000001000","000000000000001001","111111111111110000","111111111111110111","111111111111111110","000000000000010000","111111111111111100","000000000000001110","000000000000000111","000000000000001101","111111111111111110","000000000000001000","000000000000010011","000000000000001101","000000000000000010","000000000000010001","000000000000001100","000000000000010001","111111111111111101","111111111111110110","111111111111110001","000000000000000110","000000000000001011","000000000000000101","000000000000010100","000000000000010100","111111111111111001","000000000000000000","111111111111110010","000000000000000010","111111111111111100","000000000000000001","000000000000000000","000000000000000100","000000000000001010","000000000000000010","111111111111110001","000000000000000101","111111111111101100","000000000000001110","111111111111110101","111111111111110011","111111111111110111","111111111111110111","000000000000000110","111111111111110010","000000000000001000","111111111111101110","000000000000010001","111111111111110000","111111111111110101","000000000000000010","000000000000001110","111111111111110111","111111111111110011","000000000000000101","111111111111111001","000000000000010000","111111111111111010","000000000000000110","000000000000001001","000000000000001100","000000000000000110","000000000000000010","111111111111111011","000000000000000111","000000000000000001","111111111111110111","000000000000000101","111111111111110001","111111111111111000","000000000000001011","000000000000001111","111111111111110100","111111111111111000","111111111111111101","000000000000000011","111111111111110111","000000000000010011","000000000000001111","000000000000001001","000000000000001111","000000000000000000","000000000000001111","111111111111111110","000000000000000010","111111111111110100","000000000000001001","000000000000001111","000000000000010011","000000000000010000","000000000000001101","000000000000001100","000000000000010000","000000000000000111","000000000000010000","000000000000010000","111111111111101100","111111111111111100","111111111111111011","000000000000000001","111111111111110001","111111111111111000","000000000000000000","000000000000010010","000000000000000110","111111111111110110","111111111111111101","000000000000001101","000000000000010011","111111111111111111","000000000000010100"),
("111111111111111000","000000000000010011","111111111111111101","000000000000001100","000000000000010001","111111111111111101","000000000000001110","000000000000000001","111111111111111101","000000000000000000","111111111111101100","111111111111111111","111111111111101110","000000000000000000","000000000000010000","111111111111110110","111111111111111000","111111111111111101","111111111111111111","000000000000000100","111111111111110011","111111111111110001","000000000000010001","111111111111111111","111111111111110010","000000000000000101","111111111111110010","000000000000010010","000000000000001111","111111111111111100","000000000000001110","000000000000010001","111111111111111100","111111111111110001","000000000000010001","000000000000001001","000000000000000111","111111111111101101","111111111111110001","000000000000000110","111111111111111101","111111111111101110","000000000000000111","111111111111110100","000000000000001000","111111111111110100","000000000000001011","000000000000000010","111111111111101111","000000000000000110","111111111111111001","111111111111110011","111111111111110101","111111111111110100","000000000000001101","000000000000001111","111111111111110111","000000000000000110","000000000000000001","111111111111111101","000000000000001000","000000000000001010","000000000000001111","111111111111110001","000000000000000000","000000000000000011","111111111111110101","000000000000010100","000000000000001101","111111111111110111","000000000000010001","000000000000000100","000000000000001111","111111111111110111","111111111111110111","111111111111101101","111111111111111011","000000000000001000","000000000000000000","111111111111110101","000000000000001100","000000000000000010","111111111111110100","000000000000001010","000000000000000111","000000000000010011","000000000000001010","111111111111110100","000000000000000100","111111111111101111","000000000000001110","000000000000010100","000000000000001101","111111111111101100","000000000000000000","000000000000000100","111111111111111110","111111111111110111","111111111111110111","000000000000000000","111111111111111011","000000000000000000","000000000000010000","111111111111110100","111111111111101101","000000000000000010","111111111111101111","111111111111111000","000000000000000101","111111111111110101","111111111111101101","111111111111111000","000000000000000010","111111111111101100","000000000000001011","000000000000000111","111111111111110100","111111111111110110","111111111111111101","111111111111101110","111111111111110011","000000000000000000","000000000000000000","000000000000000101","111111111111110101","000000000000001101","111111111111110000","000000000000000010"),
("000000000000001110","000000000000010000","000000000000001111","111111111111110011","000000000000001010","111111111111110001","111111111111111000","000000000000000000","000000000000000111","111111111111110010","000000000000000100","000000000000010001","000000000000000000","000000000000001011","000000000000001001","111111111111111010","111111111111101100","111111111111111101","000000000000000001","000000000000010100","000000000000000000","000000000000001000","111111111111111100","111111111111110010","111111111111111101","111111111111110011","111111111111111110","111111111111111011","111111111111111010","000000000000000000","000000000000001010","000000000000001110","000000000000000001","111111111111110110","111111111111111110","111111111111111001","111111111111110011","000000000000010001","111111111111110110","000000000000001010","000000000000000010","000000000000010001","000000000000000000","000000000000010011","000000000000010011","111111111111111001","000000000000001101","000000000000000100","111111111111111001","000000000000000010","000000000000010001","000000000000000010","111111111111111110","111111111111110001","000000000000001000","000000000000000101","111111111111110011","000000000000001101","000000000000000111","111111111111110101","111111111111111110","111111111111111000","000000000000000000","111111111111111101","111111111111110100","000000000000001100","111111111111101101","111111111111111001","111111111111111011","000000000000000101","111111111111110110","000000000000001001","000000000000001001","000000000000000000","000000000000000010","000000000000010010","000000000000000101","111111111111110100","111111111111111101","111111111111101100","111111111111110000","111111111111110011","000000000000000010","111111111111111010","111111111111111101","111111111111101100","111111111111101100","111111111111111011","111111111111111001","000000000000000011","111111111111101110","111111111111110100","000000000000001010","000000000000010000","000000000000001101","000000000000001111","111111111111101101","000000000000000000","000000000000001111","000000000000010001","000000000000000110","000000000000001010","000000000000000001","111111111111110101","111111111111110111","000000000000010001","000000000000001110","111111111111101110","000000000000010000","111111111111111000","000000000000000111","000000000000001111","000000000000001111","000000000000001011","000000000000000001","000000000000000001","111111111111110010","111111111111111110","111111111111111000","000000000000000011","111111111111111110","111111111111111001","111111111111110010","000000000000000110","000000000000001111","111111111111110011","111111111111110011","000000000000000000"),
("000000000000001100","111111111111111100","000000000000001110","000000000000001111","000000000000001101","111111111111111010","111111111111110010","111111111111110011","111111111111110010","000000000000000000","000000000000000111","111111111111111101","000000000000001101","000000000000010011","111111111111101101","000000000000001110","111111111111101100","000000000000000001","000000000000010011","000000000000000001","111111111111111101","111111111111111111","111111111111110110","111111111111111010","111111111111111001","000000000000010001","111111111111111001","000000000000001010","111111111111110111","111111111111101111","000000000000000111","111111111111101110","111111111111110111","111111111111111101","111111111111111010","000000000000010011","000000000000010000","111111111111101110","000000000000001101","111111111111110100","000000000000000000","000000000000001101","000000000000000100","111111111111110110","111111111111110101","111111111111110110","111111111111110010","000000000000001000","000000000000000001","111111111111110000","111111111111110101","111111111111101110","111111111111110100","111111111111101101","000000000000001000","111111111111101111","000000000000000100","000000000000001011","000000000000010000","111111111111110011","000000000000001010","000000000000010011","111111111111101111","000000000000000000","111111111111101100","000000000000001110","000000000000000111","000000000000001010","111111111111110011","111111111111110000","111111111111111011","000000000000001101","111111111111110110","000000000000000011","111111111111110111","111111111111110000","111111111111110100","111111111111110010","000000000000001001","000000000000000010","000000000000001011","111111111111101111","000000000000000111","111111111111110000","111111111111101101","000000000000010000","111111111111111001","000000000000001111","000000000000000000","000000000000001001","111111111111110000","000000000000001100","000000000000001101","000000000000000110","000000000000001101","111111111111111000","111111111111111000","111111111111111110","111111111111110111","111111111111111001","000000000000001011","000000000000001010","000000000000001000","000000000000010001","000000000000000101","000000000000000101","000000000000000111","000000000000010100","000000000000000110","000000000000010000","000000000000000001","111111111111110111","111111111111111001","111111111111110011","000000000000001100","111111111111101110","000000000000001011","111111111111110000","111111111111111000","000000000000001000","000000000000000100","000000000000000000","000000000000010100","111111111111111110","000000000000000111","000000000000000001","111111111111111011","111111111111110000"),
("111111111111110010","111111111111110110","000000000000010100","000000000000001011","111111111111110101","000000000000001000","000000000000000001","111111111111101111","000000000000000000","000000000000000100","000000000000010000","000000000000000101","111111111111111110","000000000000001001","000000000000000001","111111111111110100","000000000000000000","000000000000000011","000000000000000100","000000000000001111","111111111111110010","111111111111111100","111111111111111011","000000000000010011","111111111111101101","000000000000000100","111111111111110001","111111111111101101","000000000000000110","111111111111111100","111111111111101101","111111111111111110","000000000000000111","111111111111111001","000000000000000100","000000000000001111","000000000000010011","111111111111110010","000000000000010100","000000000000001111","111111111111101100","000000000000000110","000000000000001101","000000000000000111","000000000000000000","111111111111110100","000000000000000101","000000000000010010","111111111111111001","111111111111101111","111111111111110110","000000000000010001","000000000000000000","000000000000001110","000000000000000110","000000000000010010","111111111111101101","000000000000010010","000000000000010100","111111111111110010","000000000000001111","000000000000010011","111111111111110111","000000000000001110","000000000000010100","111111111111110110","000000000000010010","000000000000001001","000000000000001001","000000000000000000","111111111111111010","000000000000010100","000000000000001011","000000000000001100","111111111111110010","111111111111111011","000000000000001111","111111111111110111","111111111111101100","111111111111111100","000000000000000010","000000000000010011","000000000000001101","000000000000001100","111111111111110001","111111111111101100","111111111111110101","111111111111111000","000000000000001110","111111111111111111","000000000000001101","000000000000001011","000000000000001110","000000000000001001","111111111111101101","111111111111111010","111111111111101100","111111111111111110","111111111111111011","111111111111101110","111111111111110110","111111111111110110","000000000000000000","111111111111110101","111111111111111010","000000000000010000","000000000000010001","111111111111111110","000000000000010000","111111111111110001","111111111111101111","000000000000010100","111111111111110000","111111111111111100","111111111111110111","000000000000000011","111111111111110011","111111111111110101","111111111111111001","111111111111111010","000000000000001001","000000000000000101","000000000000000110","111111111111111001","000000000000000000","111111111111111011","000000000000001110","000000000000010010"),
("000000000000000000","000000000000000011","000000000000000100","000000000000000100","000000000000001010","000000000000001111","000000000000001110","000000000000001001","111111111111110100","000000000000010010","000000000000001011","111111111111110010","111111111111111011","111111111111110001","000000000000000000","111111111111111001","000000000000000100","000000000000001011","000000000000010010","000000000000000110","111111111111111100","111111111111111111","111111111111111001","111111111111110101","111111111111111000","000000000000000000","000000000000000110","111111111111110011","000000000000000001","111111111111111110","000000000000000111","000000000000010011","000000000000000111","000000000000001101","111111111111111111","000000000000000000","000000000000000111","000000000000001011","000000000000001110","000000000000000010","111111111111111011","000000000000001010","111111111111111011","000000000000001010","111111111111110000","111111111111110100","111111111111110010","111111111111110010","111111111111101111","111111111111101101","000000000000001001","111111111111111110","000000000000010100","111111111111111010","000000000000010000","111111111111101110","111111111111111011","000000000000000101","111111111111111010","111111111111111010","000000000000010011","000000000000001111","111111111111110101","111111111111111011","000000000000000010","000000000000010010","111111111111110101","111111111111111000","111111111111110000","111111111111111100","111111111111101100","000000000000010011","000000000000000000","000000000000001111","000000000000001110","000000000000001110","111111111111110001","000000000000000000","111111111111111001","111111111111111010","000000000000010000","000000000000001100","000000000000010010","000000000000000000","111111111111111110","000000000000010100","000000000000001000","111111111111111001","111111111111111010","000000000000000011","111111111111101101","000000000000000101","000000000000001101","111111111111111101","111111111111101100","000000000000000101","111111111111110011","111111111111110010","111111111111110101","111111111111101100","111111111111111100","000000000000000001","000000000000000101","111111111111101111","000000000000001100","000000000000010001","000000000000001100","000000000000000111","000000000000000011","111111111111111111","000000000000000001","111111111111110110","000000000000000111","111111111111110110","111111111111110110","111111111111101111","000000000000000101","000000000000010001","000000000000010010","111111111111111001","000000000000010100","111111111111101100","000000000000010001","000000000000001111","000000000000001010","000000000000000000","000000000000001010","000000000000010011"),
("000000000000001001","111111111111111011","000000000000001111","111111111111111010","111111111111101111","111111111111111111","000000000000000000","000000000000001001","000000000000000000","111111111111111001","000000000000001101","000000000000010010","000000000000010001","111111111111110011","111111111111111000","000000000000000011","000000000000000110","111111111111111111","000000000000000011","111111111111111100","000000000000010010","000000000000010001","111111111111111010","111111111111110001","111111111111111100","000000000000001110","000000000000001101","111111111111110000","000000000000001011","000000000000001000","111111111111111010","111111111111111111","000000000000001011","000000000000001111","000000000000000100","111111111111110011","111111111111110101","111111111111111111","000000000000000010","000000000000000000","000000000000000000","000000000000001100","111111111111111000","111111111111110011","000000000000000100","111111111111111001","111111111111110001","000000000000000110","000000000000010100","000000000000000111","000000000000010100","111111111111111111","111111111111111010","000000000000000101","111111111111111101","000000000000001000","000000000000001111","111111111111110010","000000000000001111","000000000000001011","111111111111110000","000000000000000011","111111111111101111","000000000000000000","111111111111101101","000000000000010000","000000000000000010","000000000000001110","000000000000000001","000000000000001011","000000000000001001","111111111111111110","111111111111110000","000000000000000010","111111111111101110","000000000000001010","000000000000000110","111111111111111111","111111111111111010","111111111111111110","000000000000000001","111111111111110011","111111111111111100","111111111111110100","000000000000000111","000000000000001000","111111111111111010","000000000000010011","000000000000001010","000000000000001111","000000000000001010","111111111111101101","000000000000000111","111111111111111000","000000000000001111","111111111111101101","000000000000000111","111111111111110011","000000000000000110","000000000000000111","111111111111110001","111111111111111001","111111111111111101","000000000000001000","111111111111110001","000000000000001110","000000000000000111","111111111111101110","111111111111111111","000000000000010100","111111111111110001","111111111111111010","111111111111110110","000000000000001000","111111111111110110","111111111111110010","000000000000000110","111111111111110110","111111111111110110","111111111111110001","000000000000010011","000000000000001100","000000000000000011","000000000000000011","000000000000001001","000000000000001100","000000000000000010","000000000000010011"),
("000000000000000000","000000000000000100","000000000000000100","000000000000010100","000000000000000101","111111111111110110","000000000000010000","000000000000001101","000000000000000010","000000000000010000","111111111111101100","000000000000000010","000000000000000011","111111111111101101","111111111111101101","000000000000000111","000000000000010000","000000000000000011","000000000000001111","111111111111111100","111111111111110011","000000000000000101","111111111111111100","000000000000010010","000000000000010001","000000000000010010","111111111111101101","000000000000001101","000000000000010000","000000000000000110","000000000000000000","111111111111111000","111111111111111110","111111111111111010","111111111111110110","000000000000000000","111111111111110110","000000000000000111","000000000000001100","111111111111110011","111111111111110011","000000000000010100","000000000000000110","000000000000000000","111111111111110111","000000000000010010","000000000000000101","000000000000000010","111111111111101110","000000000000001011","000000000000000001","000000000000000111","111111111111111110","111111111111110000","000000000000010011","000000000000000010","111111111111111110","111111111111110001","000000000000001110","111111111111111110","111111111111111010","000000000000001000","111111111111110010","000000000000000001","111111111111111011","000000000000001010","000000000000000100","111111111111110101","000000000000000001","000000000000010011","111111111111111101","000000000000000101","111111111111111100","111111111111101110","111111111111110100","000000000000010011","000000000000001001","111111111111110010","000000000000000101","111111111111101100","111111111111110000","000000000000001000","000000000000001100","111111111111110011","000000000000001000","000000000000001111","000000000000001110","111111111111101111","000000000000000001","000000000000000000","000000000000000000","111111111111111001","111111111111110010","000000000000001011","000000000000000101","000000000000001100","000000000000001101","111111111111111100","111111111111110011","000000000000010001","111111111111110111","111111111111110010","000000000000010010","000000000000010010","000000000000001101","000000000000001000","000000000000000000","000000000000000100","000000000000010010","111111111111111111","111111111111110010","111111111111101111","000000000000001100","111111111111110110","111111111111111010","000000000000000101","000000000000001110","000000000000001010","111111111111110000","000000000000000000","000000000000001101","111111111111111001","000000000000010000","000000000000001111","000000000000000011","000000000000001000","111111111111110010","000000000000010001"),
("000000000000000100","111111111111111000","111111111111110100","111111111111111011","111111111111110100","111111111111111101","111111111111110010","000000000000001000","000000000000000000","000000000000010010","000000000000000011","000000000000010010","111111111111110111","000000000000001111","111111111111101100","111111111111110100","000000000000000101","000000000000001000","000000000000010011","000000000000001101","000000000000001011","111111111111111001","111111111111101110","111111111111111111","000000000000001001","111111111111111011","111111111111101101","000000000000001101","000000000000010011","111111111111101110","000000000000001100","000000000000000011","000000000000000110","111111111111101111","000000000000001000","000000000000000101","000000000000010011","000000000000010000","111111111111111010","000000000000001110","000000000000001010","000000000000001100","111111111111110100","000000000000001100","111111111111101100","000000000000001100","000000000000010000","111111111111110101","111111111111101111","111111111111111101","000000000000010001","000000000000001111","111111111111110101","111111111111111010","000000000000010000","000000000000000010","000000000000000110","000000000000010100","000000000000001000","111111111111110111","000000000000000000","000000000000001000","111111111111111110","111111111111110100","111111111111101110","111111111111101100","000000000000000000","111111111111110000","000000000000001101","000000000000000000","111111111111101111","111111111111110100","111111111111110011","000000000000010010","111111111111110110","000000000000010001","111111111111111111","111111111111111110","111111111111111000","111111111111110111","000000000000001000","111111111111101110","111111111111111000","111111111111110111","111111111111101111","111111111111110010","000000000000001000","000000000000001100","000000000000000001","000000000000000110","111111111111101110","000000000000000000","111111111111101110","111111111111111011","000000000000000000","000000000000000011","000000000000000001","111111111111111111","111111111111111010","111111111111110100","111111111111101111","000000000000000111","000000000000001010","111111111111111110","000000000000001010","000000000000010000","111111111111101101","111111111111111110","111111111111111000","111111111111110101","111111111111110000","111111111111110111","000000000000001111","111111111111110110","111111111111111100","000000000000010001","111111111111111111","000000000000010000","111111111111111111","111111111111111110","000000000000000101","111111111111111101","000000000000010000","000000000000001111","000000000000000110","111111111111101100","111111111111110111","111111111111101111"),
("000000000000000001","000000000000010011","000000000000000101","111111111111111111","111111111111110101","111111111111110110","111111111111101111","000000000000010010","000000000000001000","111111111111111111","000000000000001111","111111111111110101","000000000000010001","000000000000001110","000000000000000000","000000000000010011","000000000000000000","111111111111110001","111111111111111001","000000000000010001","111111111111110010","000000000000000110","111111111111110000","000000000000010010","000000000000001100","111111111111111001","000000000000001001","000000000000000111","000000000000001111","000000000000010011","111111111111111110","000000000000000001","111111111111111100","111111111111111100","000000000000000110","000000000000000010","000000000000001000","000000000000001001","000000000000001111","111111111111101100","000000000000001100","000000000000010000","111111111111111111","000000000000000110","000000000000010011","000000000000000001","111111111111110110","000000000000010011","000000000000001101","000000000000001100","000000000000000000","000000000000000000","000000000000010001","000000000000000100","111111111111110011","111111111111111000","000000000000000111","111111111111111111","111111111111110010","000000000000000100","000000000000000000","000000000000001000","000000000000010011","000000000000000010","000000000000001010","000000000000000100","000000000000001100","000000000000000001","111111111111110111","000000000000000101","000000000000001110","000000000000001011","111111111111110011","000000000000000000","111111111111111110","111111111111111101","111111111111110000","000000000000001001","000000000000000000","111111111111110011","000000000000001100","000000000000010001","000000000000000111","000000000000001011","000000000000000101","111111111111111101","111111111111110010","000000000000001110","000000000000000000","000000000000000011","000000000000010100","111111111111101110","111111111111110000","111111111111110010","111111111111110111","111111111111111011","111111111111111110","111111111111111110","000000000000001001","111111111111111001","000000000000010000","000000000000001101","000000000000001101","000000000000000111","000000000000010000","000000000000010011","111111111111110110","111111111111110010","000000000000001111","000000000000000011","111111111111101100","111111111111111101","111111111111110010","000000000000000011","000000000000000101","000000000000001010","000000000000001110","111111111111111001","000000000000010100","111111111111110100","111111111111101101","000000000000001101","111111111111110100","111111111111110010","111111111111110110","000000000000010100","000000000000001011","111111111111111100"),
("111111111111111010","111111111111110110","111111111111101111","111111111111110000","000000000000001110","000000000000010101","000000000000000110","111111111111101110","000000000000001101","111111111111110100","111111111111111001","000000000000000111","111111111111110001","111111111111101100","000000000000010100","000000000000001011","111111111111101011","000000000000000000","000000000000000000","111111111111101111","111111111111110100","111111111111111101","000000000000000101","000000000000000100","111111111111110010","000000000000000011","000000000000001100","111111111111110101","111111111111111111","111111111111111010","111111111111110110","000000000000010101","000000000000000100","000000000000010100","111111111111101110","000000000000001101","000000000000001101","111111111111111111","111111111111110001","111111111111110000","000000000000000110","111111111111111100","000000000000011101","000000000000001110","000000000000000000","000000000000000001","000000000000011010","111111111111111101","000000000000000110","000000000000001010","111111111111111111","111111111111110111","111111111111110001","111111111111110010","111111111111111011","000000000000000110","111111111111111011","111111111111101111","111111111111110011","111111111111110010","111111111111110000","000000000000001110","111111111111110000","111111111111111011","000000000000000011","111111111111110101","000000000000001011","111111111111111100","111111111111110001","000000000000001101","111111111111111010","000000000000000000","000000000000010001","111111111111111010","000000000000011001","000000000000010100","111111111111110011","111111111111101111","000000000000001100","000000000000000100","111111111111101111","111111111111110101","000000000000001111","111111111111110001","111111111111110010","111111111111110111","000000000000000000","111111111111111110","000000000000000100","000000000000000001","000000000000001111","000000000000000111","111111111111111010","000000000000000101","111111111111100111","000000000000000111","111111111111111001","000000000000010011","000000000000010000","111111111111110011","000000000000011000","111111111111110100","000000000000010000","000000000000000000","111111111111110110","111111111111111001","111111111111110110","000000000000010000","111111111111101010","111111111111101010","111111111111100111","000000000000001011","000000000000000100","000000000000001010","000000000000001100","111111111111110101","000000000000000101","111111111111110001","111111111111110110","111111111111111111","111111111111111101","000000000000001111","000000000000001110","000000000000000111","111111111111101110","000000000000010111","000000000000000010","111111111111111100"),
("000000000000001111","000000000000010000","111111111111011011","111111111111110111","111111111111111001","000000000000011110","000000000000010101","111111111111111000","111111111111110010","000000000000001100","000000000000010000","000000000000100010","000000000000010010","111111111111111111","000000000000100110","000000000000010000","111111111111100100","111111111111101101","000000000000001001","111111111111111010","111111111111111000","111111111111101110","111111111111110101","000000000000000100","000000000000001110","000000000000011100","111111111111111011","000000000000000011","111111111111111001","000000000000000101","111111111111111010","000000000000010001","111111111111110001","111111111111110000","000000000000010100","000000000000000100","111111111111110111","111111111111101100","000000000000000111","000000000000000101","111111111111110110","000000000000000011","000000000000001000","000000000000000101","111111111111101100","111111111111101110","111111111111111110","000000000000001110","111111111111110010","111111111111110111","000000000000001010","111111111111110010","000000000000001000","111111111111100111","000000000000000000","111111111111011110","000000000000000010","111111111111110011","111111111111111011","000000000000000010","111111111111111101","111111111111111010","111111111111111010","111111111111101101","000000000000001111","111111111111110000","111111111111111100","000000000000011011","111111111111110111","000000000000000110","000000000000000000","000000000000010000","111111111111110101","111111111111111110","000000000000010000","000000000000011010","111111111111110000","000000000000001011","111111111111100101","111111111111011110","111111111111111111","111111111111111000","111111111111011100","111111111111111110","000000000000000110","000000000000000000","111111111111100001","000000000000001111","000000000000000100","000000000000001100","000000000000011010","111111111111111011","000000000000100001","111111111111111111","111111111111111100","111111111111111101","111111111111110110","000000000000010001","111111111111110110","111111111111100011","000000000000010100","000000000000000100","000000000000000010","111111111111111001","111111111111110100","111111111111111010","000000000000000101","000000000000010101","000000000000000010","111111111111100101","000000000000000000","111111111111110101","000000000000001111","111111111111110111","111111111111100011","000000000000011110","000000000000010101","000000000000000100","000000000000000000","000000000000001100","000000000000001111","111111111111111000","000000000000011101","000000000000001011","000000000000000000","000000000000011110","000000000000010110","111111111111011110"),
("000000000000010100","000000000000011001","111111111111110110","000000000000010110","111111111111011110","000000000000001101","000000000000001010","111111111111101100","000000000000001001","000000000000001001","111111111111110101","000000000000000000","000000000000010011","000000000000010000","000000000000000001","111111111111111111","111111111111011101","111111111111101101","000000000000000000","000000000000000101","111111111111110011","111111111111111000","111111111111100111","000000000000000000","000000000000000001","111111111111111110","111111111111110110","000000000000010000","111111111111111011","000000000000010111","111111111111110101","000000000000000010","111111111111111111","000000000000010000","000000000000001111","111111111111101100","000000000000001001","000000000000000000","000000000000000110","111111111111101110","000000000000010000","000000000000001111","000000000000010101","000000000000010101","111111111111111011","111111111111110011","000000000000100100","000000000000100111","000000000000000001","000000000000010111","000000000000000011","000000000000000000","000000000000000010","111111111111100000","000000000000000110","111111111111011110","111111111111101111","111111111111111010","111111111111101101","111111111111110010","111111111111110100","111111111111101111","111111111111110000","000000000000000011","000000000000000101","111111111111110000","111111111111110101","000000000000100010","111111111111101001","000000000000000110","000000000000000001","000000000000001011","111111111111101000","111111111111100010","000000000000011000","000000000000000001","111111111111100010","111111111111111010","111111111111111110","111111111111100011","111111111111101101","111111111111100001","111111111111110101","111111111111111111","111111111111100111","111111111111111000","111111111111100111","000000000000000000","000000000000001101","111111111111110101","000000000000011100","000000000000010011","000000000000010101","000000000000001000","111111111111011010","000000000000000010","111111111111111011","000000000000000000","000000000000000101","111111111111101111","000000000000010000","000000000000000010","111111111111111011","000000000000000101","000000000000001000","111111111111111111","111111111111111001","000000000000100101","111111111111111001","111111111111011100","111111111111101110","111111111111111110","000000000000011100","111111111111111101","111111111111110110","000000000000100010","000000000000000110","111111111111101011","111111111111110000","000000000000000001","111111111111110100","000000000000000001","000000000000001100","000000000000010000","000000000000100100","000000000000010111","111111111111110011","111111111111101110"),
("111111111111110000","000000000000011011","111111111111110000","111111111111111101","111111111111111000","000000000000010110","000000000000011110","111111111111111011","111111111111111011","111111111111111111","000000000000001000","000000000000000011","000000000000001111","111111111111100111","000000000000000010","111111111111110101","111111111111110111","000000000000010000","000000000000001100","111111111111110101","111111111111110110","000000000000010100","000000000000000100","000000000000000101","000000000000010101","111111111111111100","000000000000000110","000000000000000000","111111111111100101","000000000000000001","111111111111110101","000000000000100001","111111111111111010","000000000000011110","000000000000010110","111111111111111101","000000000000000000","000000000000010000","111111111111111001","111111111111101001","111111111111110110","000000000000000001","000000000000001101","000000000000011010","111111111111100000","000000000000000110","000000000000010101","000000000000000101","111111111111101111","000000000000001110","111111111111110101","000000000000000110","000000000000001011","000000000000000000","111111111111110111","111111111111100000","000000000000010000","111111111111110001","111111111111111110","111111111111111100","111111111111110100","000000000000000100","000000000000001011","111111111111111101","000000000000001011","000000000000001001","000000000000001000","000000000000011000","000000000000000110","111111111111111111","000000000000001110","111111111111111100","111111111111111101","111111111111100100","000000000000011011","111111111111111101","111111111111110100","000000000000000000","111111111111110000","111111111111101000","111111111111101101","000000000000000000","000000000000000001","000000000000000001","111111111111111011","111111111111100001","000000000000000001","000000000000010000","000000000000000011","111111111111110010","000000000000010100","000000000000100101","000000000000001000","000000000000000101","000000000000000011","000000000000010000","000000000000010011","000000000000001000","000000000000011001","000000000000000000","000000000000000001","000000000000000000","000000000000010010","111111111111111001","111111111111110101","111111111111111101","111111111111100101","000000000000000011","111111111111111100","111111111111101110","000000000000000000","000000000000000100","000000000000011111","000000000000001010","111111111111011110","000000000000000111","000000000000001111","111111111111111110","111111111111101010","111111111111111100","000000000000000001","000000000000000111","000000000000010001","000000000000100011","000000000000000100","000000000000000011","000000000000000001","111111111111101010"),
("111111111111110111","000000000000001001","111111111111011010","111111111111111101","000000000000001011","000000000000001111","000000000000000100","111111111111111101","111111111111111000","000000000000011000","111111111111111111","000000000000010110","000000000000001110","111111111111111010","000000000000001101","000000000000010100","111111111111111100","000000000000001011","000000000000000000","000000000000000111","111111111111110010","111111111111111010","111111111111110000","111111111111110100","000000000000000001","000000000000000011","111111111111110110","000000000000010011","000000000000001000","111111111111110100","111111111111100100","000000000000000010","000000000000000001","000000000000011011","000000000000010010","000000000000001000","111111111111111001","111111111111111011","111111111111110011","111111111111111100","111111111111110001","000000000000010000","000000000000010100","000000000000100011","111111111111111111","111111111111110001","000000000000001110","000000000000010010","111111111111101000","000000000000011010","111111111111110010","000000000000000001","111111111111111111","111111111111110011","111111111111111110","111111111111011111","111111111111101001","111111111111110001","111111111111101100","111111111111111110","000000000000000011","000000000000000110","111111111111111101","111111111111101000","111111111111110011","111111111111110001","111111111111110001","000000000000010100","111111111111110001","111111111111101100","000000000000010011","111111111111110100","111111111111110011","111111111111100111","000000000000010011","000000000000011011","000000000000000010","000000000000010111","111111111111111010","111111111111101010","000000000000000101","111111111111100110","111111111111110111","000000000000000101","000000000000000000","111111111111111011","111111111111111110","000000000000000011","000000000000001111","000000000000010010","111111111111110110","000000000000010001","000000000000010011","000000000000010010","111111111111011111","111111111111110110","000000000000000011","000000000000100101","000000000000001100","111111111111101000","000000000000010011","000000000000010100","000000000000010001","000000000000001100","000000000000010001","000000000000000101","111111111111110000","000000000000010001","111111111111111001","111111111111110110","111111111111101011","111111111111111111","000000000000011001","111111111111111001","111111111111011110","000000000000100000","000000000000001101","000000000000000010","000000000000001011","111111111111111100","000000000000011010","000000000000000000","111111111111111100","000000000000010011","000000000000000000","000000000000010011","000000000000011010","111111111111101101"),
("000000000000011000","000000000000110110","111111111111111011","111111111111111101","000000000000011011","111111111111110011","000000000000001011","111111111111100110","000000000000001001","000000000000000100","000000000000000000","000000000000101110","111111111111110101","000000000000001011","000000000000110010","000000000000001100","111111111111101111","111111111111101101","111111111111110101","111111111111110110","000000000000001010","111111111111101111","111111111111110001","111111111111110010","000000000000000010","000000000000000101","000000000000000001","000000000000010000","111111111111110010","000000000000010100","111111111111010101","000000000000000001","111111111111100100","000000000000000011","111111111111111101","000000000000000111","000000000000011011","111111111111100001","111111111111110100","111111111111011111","000000000000001100","000000000000011100","000000000000011100","111111111111111100","111111111111110101","000000000000000001","000000000000010111","000000000000100000","111111111111110100","000000000000001111","000000000000000110","111111111111110010","000000000000001001","111111111111111001","000000000000000110","111111111111100000","000000000000000010","000000000000000010","111111111111101111","000000000000010000","000000000000001100","000000000000000110","111111111111110110","111111111111101111","111111111111101001","000000000000001001","111111111111110100","000000000000011110","111111111111001101","111111111111101010","000000000000100000","111111111111110001","000000000000000111","111111111111011011","000000000000100000","111111111111111111","111111111111110111","111111111111111110","000000000000000010","111111111111111001","000000000000001100","111111111111111110","000000000000001001","111111111111111111","000000000000000000","000000000000001010","111111111111101010","000000000000000101","000000000000011011","111111111111111000","111111111111111110","000000000000000001","000000000000011001","111111111111111001","111111111111110001","000000000000011001","111111111111111111","000000000000000100","000000000000010110","000000000000000011","000000000000011011","000000000000010100","111111111111111110","111111111111101011","111111111111110010","111111111111111111","111111111111100100","000000000000010100","111111111111100101","111111111111110111","111111111111101010","111111111111110101","000000000000010000","111111111111101100","111111111111011110","000000000000001001","000000000000011000","111111111111101001","000000000000001000","111111111111100100","000000000000000001","111111111111011011","000000000000010011","000000000000011010","111111111111110001","000000000000001111","000000000000001001","111111111111101111"),
("000000000000011011","000000000000010010","111111111111111110","111111111111111110","000000000000011101","000000000000010100","000000000000001001","111111111111100111","000000000000000110","000000000000001011","111111111111101100","000000000000001010","000000000000000100","000000000000001000","000000000000000100","000000000000010100","111111111111101110","111111111111111001","111111111111111100","111111111111110011","111111111111101011","111111111111111111","000000000000001100","000000000000000100","000000000000011000","000000000000001000","111111111111111101","111111111111111010","111111111111111001","111111111111111010","111111111111101011","000000000000000111","111111111111101011","000000000000000111","111111111111111111","111111111111101110","000000000000001101","111111111111111011","111111111111100011","000000000000000000","111111111111111010","000000000000000010","000000000000110001","000000000000001000","111111111111110000","111111111111100010","000000000000011011","000000000000011011","111111111111110000","000000000000011100","000000000000011001","111111111111101101","000000000000001110","000000000000001000","111111111111110111","111111111111011010","111111111111110011","111111111111101100","000000000000000000","111111111111111100","000000000000001101","111111111111011111","111111111111111111","111111111111111111","000000000000001111","000000000000001000","000000000000001110","000000000000001111","111111111111001011","000000000000010000","000000000000000110","000000000000000001","000000000000011001","111111111111101100","111111111111111101","000000000000011011","111111111111011110","000000000000000110","111111111111100110","111111111111111101","000000000000010001","111111111111111001","000000000000010011","000000000000000001","111111111111110000","000000000000000111","111111111111101100","000000000000001010","000000000000010101","000000000000010110","000000000000000100","000000000000000101","000000000000010000","000000000000100000","111111111111110110","111111111111111010","000000000000001000","111111111111110110","000000000000000001","111111111111100110","111111111111111110","000000000000010100","000000000000000100","000000000000000001","111111111111110100","000000000000100110","111111111111011101","000000000000001110","111111111111111010","000000000000000111","000000000000000100","111111111111100011","000000000000000100","000000000000000101","111111111111010100","000000000000001011","000000000000100001","111111111111101011","000000000000000011","000000000000000001","000000000000001000","000000000000000100","000000000000000101","000000000000000010","000000000000001100","000000000000000010","000000000000000011","111111111111110001"),
("000000000000001010","000000000000011101","111111111111110010","000000000000000010","111111111111110010","111111111111110101","000000000000010001","111111111111011010","111111111111100110","000000000000011110","000000000000000110","000000000000101111","000000000000000011","111111111111111111","000000000000000010","111111111111111110","111111111111110000","000000000000000100","000000000000010010","111111111111111011","000000000000000001","000000000000000000","000000000000010010","111111111111110001","000000000000000010","111111111111110001","111111111111101101","111111111111110101","000000000000000000","000000000000011011","111111111111011011","000000000000011100","111111111111111000","000000000000100100","111111111111100111","000000000000000111","111111111111110100","000000000000000101","111111111111111110","111111111111110111","000000000000001101","000000000000001000","000000000000010001","000000000000100101","111111111111010100","111111111111100011","000000000000001011","000000000000000111","111111111111110000","000000000000001000","111111111111110110","111111111111101010","000000000000010111","000000000000000001","111111111111011010","111111111111110110","000000000000000000","111111111111110000","111111111111110110","000000000000000011","000000000000001111","111111111111111010","111111111111110010","000000000000000110","111111111111110000","000000000000000000","000000000000000011","000000000000001001","111111111111011001","111111111111111111","000000000000011001","000000000000001000","000000000000011110","111111111111100000","000000000000011100","000000000000010001","111111111111010101","111111111111110011","111111111111111111","111111111111110110","000000000000011000","111111111111111110","000000000000000100","111111111111101010","111111111111111001","111111111111110000","111111111111110011","000000000000001101","111111111111111011","000000000000011100","000000000000000100","000000000000011110","000000000000011111","000000000000100100","111111111111100110","000000000000011110","000000000000001110","000000000000010010","111111111111111001","111111111111101010","000000000000011101","000000000000110011","000000000000001010","111111111111111100","000000000000001110","000000000000011100","111111111111101001","000000000000010001","111111111111111011","000000000000001111","111111111111110100","111111111111111111","000000000000011110","111111111111100011","111111111111100110","000000000000100000","000000000000000110","111111111111111101","111111111111101001","000000000000000011","000000000000000011","111111111111110010","000000000000010011","111111111111110001","000000000000000000","000000000000100000","000000000000000111","111111111111011111"),
("000000000000001100","000000000000011111","111111111111011001","111111111111110011","111111111111111111","111111111111111000","000000000000101010","111111111111011110","111111111111110011","000000000000101000","111111111111111111","000000000000110010","111111111111110101","111111111111100111","111111111111111111","000000000000001011","000000000000000001","000000000000001110","111111111111110111","111111111111101011","000000000000000100","000000000000100000","000000000000000100","111111111111111001","000000000000001100","000000000000001000","111111111111100011","000000000000001111","111111111111101100","000000000000010110","111111111111100001","000000000000000000","000000000000000010","000000000000100010","111111111111111000","111111111111111011","000000000000001010","111111111111011111","111111111111111000","111111111111011101","000000000000010010","111111111111111000","000000000000101110","000000000000100010","111111111111100011","111111111111011100","000000000000101011","000000000000010000","111111111111010011","000000000000011001","000000000000001000","000000000000000000","000000000000001100","111111111111100110","111111111111111101","111111111111010011","111111111111110000","000000000000001011","111111111111101110","000000000000000001","111111111111111011","000000000000000101","111111111111110100","111111111111110111","000000000000000011","000000000000010010","111111111111111010","000000000000011010","111111111111011011","111111111111110000","000000000000000100","000000000000001001","000000000000000100","111111111111011010","000000000000001001","000000000000001010","111111111111111000","000000000000001011","111111111111111000","111111111111110010","000000000000001010","111111111111111001","111111111111111000","111111111111110000","111111111111101110","111111111111111001","111111111111111000","111111111111110100","000000000000011111","000000000000001011","111111111111111011","111111111111111010","111111111111111110","000000000000011101","111111111111011000","000000000000000001","000000000000000110","000000000000001110","111111111111111111","111111111111110111","000000000000100001","000000000000010011","000000000000001011","111111111111101100","000000000000000010","000000000000100110","111111111111101110","000000000000000110","000000000000000011","000000000000001010","111111111111100111","000000000000001101","000000000000100010","111111111111010101","111111111111101100","000000000000001100","000000000000010110","111111111111101011","000000000000001101","111111111111110110","000000000000001010","111111111111111000","000000000000010101","111111111111101100","000000000000001110","000000000000100100","000000000000101111","111111111111101010"),
("111111111111100111","000000000000101010","111111111111101111","000000000000001100","111111111111101001","111111111111111101","111111111111111000","111111111111101100","000000000000001010","111111111111111101","000000000000000110","000000000000100000","000000000000001001","000000000000010000","111111111111101111","111111111111111011","111111111111110101","000000000000000000","111111111111100101","111111111111100110","000000000000001010","000000000000100110","000000000000011001","111111111111111011","000000000000001001","000000000000001011","000000000000000001","000000000000000001","000000000000001010","000000000000001110","111111111111111010","111111111111110001","111111111111111100","000000000000100001","000000000000100010","000000000000000100","111111111111101011","111111111111110101","000000000000011111","111111111111100000","111111111111111011","000000000000000001","000000000000001010","000000000000110000","000000000000001001","000000000000011000","000000000000000101","111111111111111101","111111111111110111","000000000000001010","111111111111110000","000000000000000111","111111111111110100","000000000000001101","111111111111111001","000000000000000101","000000000000001001","000000000000001010","111111111111111101","000000000000000100","111111111111100000","000000000000010110","000000000000011011","111111111111111110","000000000000001111","000000000000001111","000000000000010000","111111111111110010","111111111111111010","000000000000000000","111111111111111101","000000000000000100","111111111111100111","111111111111100110","000000000000001111","111111111111111100","111111111111111110","000000000000000111","000000000000010110","000000000000000111","111111111111101011","111111111111110100","000000000000000101","111111111111110000","000000000000100100","000000000000000011","000000000000000101","000000000000001011","000000000000001000","000000000000010100","000000000000001111","111111111111111111","111111111111011111","000000000000011111","111111111111100101","000000000000001110","000000000000000000","111111111111111000","111111111111110100","000000000000010110","111111111111101000","000000000000000001","111111111111111100","000000000000001111","000000000000100110","111111111111110100","000000000000000001","111111111111011101","111111111111011101","000000000000000100","000000000000001011","000000000000011111","111111111111011111","111111111111100000","000000000000001100","111111111111101100","111111111111101011","111111111111110101","111111111111111101","111111111111011101","000000000000001101","000000000000011110","000000000000000110","000000000000110101","000000000000000001","111111111111110111","000000000000001010","111111111111110111"),
("111111111111100100","000000000000110101","111111111111011000","000000000000010110","111111111111101001","111111111111110100","111111111111111000","000000000000000100","000000000000001111","000000000000010000","000000000000001010","000000000000001000","000000000000000010","111111111111110010","000000000000000101","000000000000011001","111111111111111111","000000000000001110","111111111111110101","111111111111100011","000000000000000111","111111111111111010","111111111110101010","000000000000001000","111111111111101111","000000000000010111","111111111111011110","111111111111110010","000000000000000000","111111111111111110","111111111111101111","000000000000010011","111111111111100110","000000000000101001","000000000000000000","111111111111111100","111111111111101001","000000000000010110","111111111111111000","111111111111010010","000000000000010110","111111111111110111","000000000000110011","000000000000100111","111111111111001110","000000000000000111","000000000000011111","000000000000011001","111111111111101111","111111111111111100","000000000000001110","111111111111100100","000000000000010110","000000000000001110","111111111111111010","111111111111010011","000000000000001100","000000000000001101","000000000000000101","000000000000010100","111111111111111111","111111111111111010","111111111111111000","111111111111111101","111111111111111111","000000000000000011","000000000000100001","000000000000000110","111111111111111111","111111111111111010","000000000000100000","000000000000011101","000000000000001001","111111111111111101","000000000000011001","111111111111110100","111111111111101010","000000000000001011","111111111111100110","111111111111110000","111111111111110010","111111111111110011","111111111111111010","111111111111110011","000000000000101000","000000000000000000","000000000000000110","111111111111111110","111111111111101111","000000000000010101","000000000000000001","000000000000001100","000000000000011101","000000000000100000","111111111111101011","111111111111101110","000000000000000101","111111111111101101","000000000000011101","111111111111111101","111111111111110000","111111111111110011","111111111111101100","000000000000001100","000000000000110001","000000000000000000","111111111111101001","111111111111110010","111111111111101101","111111111111101110","111111111111101111","111111111111101111","111111111111110001","111111111111010011","111111111111101100","111111111111111111","000000000000000010","111111111111110010","111111111111101011","111111111111101010","000000000000001010","000000000000010000","111111111111111111","000000000000110100","111111111111101111","000000000000110000","111111111111111011","111111111111011110"),
("111111111111110001","000000000000001110","111111111111100011","000000000000010111","111111111111001011","111111111111100101","000000000000100011","111111111111110111","000000000000001010","000000000000010000","000000000000000011","000000000000001011","000000000000001110","111111111111000110","111111111111100011","000000000000101001","000000000000000001","000000000000010011","000000000000011100","000000000000000111","000000000000001111","111111111111110001","111111111110110001","111111111111111100","000000000000011000","111111111111111110","111111111111110100","000000000000001010","111111111111011110","000000000000001001","000000000000000000","111111111111101000","000000000000101000","000000000000101110","111111111111110111","111111111111101011","000000000000010000","111111111111111110","111111111111110100","111111111111100000","111111111111110110","111111111111101001","000000000000110100","000000000000101110","111111111111100110","111111111111010101","000000000000011100","000000000000000111","111111111111101010","111111111111011101","000000000000000010","000000000000001111","000000000000000011","111111111111101110","000000000000000111","111111111111101111","111111111111111001","000000000000001001","111111111111110101","111111111111110000","000000000000010101","000000000000100010","000000000000011011","111111111111110110","111111111111111000","111111111111111001","111111111111101100","000000000000010011","000000000000101001","000000000000001010","000000000000001010","000000000000000010","111111111111111110","000000000000011111","111111111111101011","000000000000000110","111111111111100110","000000000000100010","111111111111011101","000000000000001010","000000000000000101","111111111111110001","000000000000010010","111111111111100000","000000000000000010","111111111111111000","111111111111101001","000000000000000000","000000000000000000","000000000000010000","111111111111111101","000000000000010010","000000000000000111","000000000000101101","111111111111100111","000000000000000001","111111111111110111","000000000000000110","111111111111111101","111111111111100101","000000000000100001","000000000000001011","000000000000010000","000000000000001110","000000000000000000","000000000000111000","111111111111010000","000000000000000010","111111111111010110","000000000000001001","111111111111010001","111111111111101101","000000000000010100","111111111111110010","111111111111010101","000000000000011010","000000000000101010","000000000000001001","111111111111110010","111111111111111000","000000000000000011","000000000000010111","000000000000001110","000000000000011010","000000000000100000","000000000000101101","000000000000011011","111111111111100001"),
("111111111111100101","000000000000001111","111111111111101101","000000000000001011","111111111111100011","111111111111110111","000000000000111001","111111111111101111","111111111111111000","000000000000101000","000000000000000110","000000000000010001","111111111111110101","111111111111010011","111111111111100111","000000000000010110","000000000000011001","000000000000000111","000000000000010001","000000000000011001","111111111111110111","111111111111101011","111111111110101111","000000000000001000","000000000000000111","000000000000001101","111111111111111000","000000000000100010","000000000000000000","111111111111111110","000000000000000000","000000000000000001","000000000000010111","000000000000100111","111111111111110010","111111111111110100","111111111111111001","111111111111110101","111111111111111101","111111111111111010","111111111111101000","000000000000000101","000000000000100110","000000000000010100","111111111111100100","111111111111100110","000000000000100011","000000000000010100","111111111111100100","111111111111011001","000000000000010110","111111111111111010","000000000000010001","000000000000000001","111111111111100110","111111111111100011","111111111111110100","000000000000010110","000000000000000100","111111111111111110","000000000000000100","000000000000001001","000000000000001110","111111111111110110","000000000000000000","111111111111110011","000000000000000000","000000000000001000","000000000000001011","111111111111110010","111111111111111111","000000000000001011","000000000000010000","111111111111111011","000000000000000111","111111111111111111","000000000000000101","000000000000100101","111111111111011100","111111111111110000","000000000000000000","000000000000000000","000000000000000111","111111111111011010","000000000000001000","000000000000000000","000000000000010001","000000000000010001","111111111111110010","111111111111110100","111111111111110111","000000000000000001","000000000000100101","000000000000101111","111111111111011110","111111111111111111","111111111111110111","111111111111111110","000000000000010111","111111111111110101","000000000000011010","111111111111110110","000000000000010111","000000000000001110","000000000000000011","000000000000100011","111111111111010111","000000000000011001","111111111111111011","000000000000010101","111111111111110100","000000000000000011","111111111111111111","111111111111100001","111111111111101011","000000000000011011","000000000000101100","000000000000000011","111111111111101110","111111111111111010","000000000000000100","000000000000100011","000000000000011011","000000000000100010","000000000000101000","000000000000101001","000000000000001100","111111111111110000"),
("000000000000100011","000000000000101100","111111111111111111","111111111111101100","111111111111101010","000000000000010001","000000000000001101","000000000000010011","111111111111011101","000000000000000111","111111111111111001","000000000000011101","111111111111110000","111111111111111011","000000000000000110","000000000000001110","111111111111100011","000000000000000110","000000000000000000","111111111111110011","111111111111111010","111111111111100110","111111111111001010","111111111111101010","000000000000011010","111111111111111011","000000000000000000","000000000000000000","111111111111111000","000000000000011100","111111111111101110","000000000000011011","111111111111010010","000000000000110011","111111111111011100","000000000000000001","111111111111110011","111111111111110100","111111111111110011","111111111111111010","111111111111111101","000000000000100010","000000000000001011","000000000000011100","111111111111100100","000000000000010010","000000000000011010","000000000000100000","111111111111110001","000000000000010101","111111111111101111","111111111111110110","000000000000110011","000000000000000001","111111111111101101","111111111111110100","000000000000100110","111111111111111111","111111111111111001","111111111111111010","000000000000100001","111111111111010101","111111111111011011","111111111111101110","111111111111110111","000000000000001000","111111111111110110","000000000000001001","111111111111011110","111111111111100111","000000000000100011","111111111111111100","000000000000110011","111111111111110000","000000000000101001","000000000000001110","111111111111101011","111111111111011011","000000000000001010","111111111111001000","000000000000001011","111111111111101101","111111111111111110","000000000000000110","111111111111111101","000000000000001000","111111111111101101","000000000000010001","000000000000001110","000000000000010111","000000000000001101","000000000000001000","000000000000011110","000000000000100101","111111111111100111","000000000000011011","000000000000001001","111111111111111100","000000000000010010","000000000000011100","000000000000010000","000000000000011000","000000000000011001","111111111111111001","000000000000001001","111111111111111101","111111111111010111","000000000000101100","000000000000000111","111111111111111101","111111111111011000","111111111111100111","000000000000100011","111111111111110011","111111111111011000","000000000000100000","000000000000100101","111111111111111010","000000000000001101","111111111111101110","000000000000001001","111111111111101111","000000000000000011","000000000000000110","111111111111111110","000000000000110010","111111111111110100","111111111111100100"),
("000000000000100000","000000000000100111","111111111111101000","111111111111110100","000000000000000010","000000000000100100","000000000000000110","111111111111101110","111111111111100100","000000000000010110","111111111111100110","000000000000000011","000000000000000000","000000000000010000","000000000000100000","000000000000001100","111111111111011010","000000000000000000","111111111111101111","111111111111010111","111111111111110100","000000000000001001","111111111111011100","111111111111110010","111111111111110010","000000000000010001","111111111111110011","111111111111101111","000000000000010111","000000000000100010","111111111111100000","000000000000100110","111111111111101101","000000000000100011","111111111111100110","000000000000001011","000000000000000001","111111111111010000","000000000000001010","111111111111101010","000000000000000101","000000000000110001","000000000000010011","000000000000000111","111111111111010110","111111111111110001","000000000000100111","000000000000100010","111111111111110011","000000000000011011","111111111111101000","111111111111011011","000000000000100011","000000000000000111","111111111111010100","111111111111011111","000000000000010000","111111111111110111","111111111111110110","000000000000000100","000000000000001101","111111111111101111","111111111111010100","111111111111110000","000000000000001010","000000000000000010","000000000000001001","000000000000011010","111111111111100011","000000000000000000","000000000000101100","111111111111101100","000000000000100010","000000000000000000","000000000000110011","000000000000011100","111111111111010011","111111111111101100","111111111111101011","111111111111001100","000000000000000000","111111111111011001","111111111111011101","000000000000000010","000000000000000101","111111111111101110","111111111111101100","000000000000000000","000000000000101100","111111111111110111","000000000000100111","000000000000010001","000000000000011101","000000000000000100","111111111111110100","000000000000001011","111111111111110101","000000000000001001","000000000000100101","000000000000001110","000000000000010000","000000000000001011","000000000000010111","111111111111110110","111111111111111001","000000000000001000","111111111111010100","000000000000110100","111111111111101100","111111111111111010","111111111111101000","111111111111101001","000000000000100111","111111111111100011","111111111111111000","000000000000001000","000000000000100011","111111111111101110","111111111111110000","111111111111101101","000000000000010101","111111111111010001","000000000000100110","000000000000010101","000000000000001101","000000000000001110","111111111111110111","111111111111011101"),
("000000000000100110","000000000000001011","111111111111010011","111111111111110011","111111111111100100","000000000000010000","000000000000010110","111111111111110001","111111111111011000","000000000000000111","111111111111101101","000000000000010010","111111111111111101","000000000000010111","000000000000010110","000000000000010101","111111111111100111","000000000000001001","000000000000001001","111111111111111000","111111111111011011","000000000000001011","111111111111111000","111111111111101110","000000000000001111","000000000000000000","000000000000000001","000000000000000000","000000000000001101","000000000000001011","111111111111111110","000000000000010000","111111111111101010","000000000000101011","111111111111101110","000000000000000000","111111111111111010","111111111111001010","111111111111111001","111111111111110100","111111111111111010","000000000000010110","000000000000001110","000000000000011101","111111111111101111","111111111111110011","000000000000001100","000000000000011100","111111111111101011","000000000000111111","111111111111110000","111111111111110011","000000000000001110","111111111111110011","111111111111011101","111111111111110001","000000000000010101","111111111111101111","111111111111101111","111111111111101101","000000000000100111","111111111111101001","111111111111010011","111111111111101100","111111111111111101","111111111111110000","000000000000100100","000000000000010001","111111111111011111","111111111111110001","000000000000011110","000000000000001011","000000000000110011","111111111111110111","000000000000011101","111111111111111100","111111111111100100","111111111111100101","000000000000000100","111111111111100110","111111111111110001","111111111111011110","111111111111101110","000000000000000101","111111111111110010","111111111111111010","111111111111110001","000000000000000110","000000000000100011","000000000000000110","000000000000000000","000000000000011011","000000000000100101","000000000000010001","111111111111010001","000000000000001100","000000000000001100","000000000000100011","000000000000010000","111111111111110000","000000000000001110","000000000000011100","000000000000011001","111111111111100110","000000000000000001","000000000000100100","111111111111110000","000000000000111101","111111111111110000","111111111111111010","111111111111010100","000000000000000110","000000000000100000","111111111111011110","111111111111001100","000000000000011000","000000000000010111","000000000000010000","111111111111110111","111111111111111011","000000000000000000","111111111111101011","000000000000100010","000000000000001110","000000000000010110","000000000000011010","111111111111111101","111111111111110111"),
("000000000000010000","000000000000001000","111111111111111011","111111111111111010","111111111111110000","000000000000100101","000000000000011010","000000000000000011","111111111111100100","000000000000001111","111111111111100111","000000000000000111","111111111111100110","000000000000100100","000000000000100111","111111111111111011","111111111111110100","000000000000000000","111111111111111101","111111111111110001","111111111111110010","000000000000000000","111111111111100001","111111111111110001","111111111111110100","000000000000011111","111111111111101011","111111111111111001","000000000000000010","000000000000000111","111111111111100001","000000000000010000","111111111111001101","000000000000100010","111111111111111101","000000000000000000","000000000000000000","111111111111110110","111111111111110101","111111111111100111","000000000000010001","000000000000010111","000000000000100010","000000000000010001","111111111111101001","111111111111111000","000000000000011010","000000000000010010","111111111111010101","000000000000010000","111111111111000111","111111111111101101","000000000000001111","000000000000000110","111111111111101101","111111111111110010","111111111111111001","000000000000000101","111111111111011001","111111111111111100","000000000000100111","111111111111101110","111111111111100100","111111111111110111","111111111111110100","000000000000000111","000000000000010010","000000000000011011","111111111111011010","111111111111100111","000000000000011010","111111111111110110","000000000000010111","111111111111110001","000000000000000010","000000000000000100","111111111111010101","000000000000000000","111111111111111100","111111111111111001","000000000000001101","111111111111110111","111111111111110000","111111111111110100","111111111111111001","000000000000000011","111111111111110110","000000000000001111","000000000000001100","000000000000001101","000000000000010000","000000000000001100","000000000000100101","000000000000010100","111111111111100111","111111111111110101","000000000000001000","000000000000011001","000000000000011001","111111111111111110","000000000000011000","000000000000100111","000000000000101001","111111111111101111","111111111111110001","000000000000010101","111111111111111000","000000000000001101","111111111111101101","111111111111101110","111111111111111000","111111111111111111","000000000000100011","111111111111101000","111111111111010001","000000000000010011","000000000000011111","000000000000001000","000000000000000011","000000000000001001","111111111111111000","111111111111010011","000000000000010100","000000000000000010","111111111111111000","000000000000011111","000000000000001111","111111111111110001"),
("000000000000011011","000000000000100101","111111111111110110","111111111111111001","000000000000000000","000000000000101010","000000000000001100","111111111111110100","111111111111111101","000000000000010110","111111111111111001","000000000000011110","000000000000001110","000000000000011100","000000000000010100","000000000000011001","111111111111110100","000000000000010000","000000000000000000","111111111111101100","000000000000000000","111111111111111000","111111111111101001","111111111111011111","111111111111111010","000000000000100000","111111111111111010","000000000000010010","000000000000001101","000000000000010100","111111111111110101","000000000000101001","111111111111110000","000000000000100010","111111111111100010","111111111111110011","000000000000010100","111111111111111011","111111111111111001","000000000000000101","111111111111111000","000000000000011010","000000000000011101","000000000000010011","111111111111011011","000000000000010001","000000000000011111","000000000000010111","111111111111011111","000000000000010110","000000000000000011","111111111111011111","000000000000011001","111111111111111001","111111111111111101","111111111111100101","000000000000000000","000000000000001011","111111111111011010","000000000000001011","000000000000100010","111111111111110000","111111111111100110","111111111111110010","111111111111110110","111111111111110100","000000000000001000","000000000000010111","111111111111110100","000000000000000101","000000000000001111","111111111111111011","000000000000101100","111111111111100011","000000000000001010","000000000000000101","111111111111011001","111111111111111110","111111111111111110","111111111111101000","111111111111110100","111111111111011110","111111111111101010","111111111111100010","111111111111101101","111111111111100110","111111111111110010","000000000000001001","000000000000100100","111111111111111001","000000000000011010","111111111111110010","000000000000011000","000000000000100100","111111111111100100","000000000000001100","000000000000001000","000000000000011010","000000000000011010","111111111111101010","000000000000000000","000000000000011000","000000000000001110","111111111111101000","111111111111110011","000000000000001110","111111111111111110","000000000000001011","111111111111101011","111111111111100000","111111111111101001","000000000000000010","000000000000001011","111111111111111111","111111111111100010","000000000000000010","000000000000011011","000000000000000001","000000000000000100","000000000000000000","111111111111111001","111111111111010110","000000000000000000","111111111111111011","000000000000011100","000000000000011010","000000000000011011","111111111111100001"),
("111111111111111110","000000000000010100","000000000000000000","000000000000000101","111111111111110100","111111111111111011","000000000000011101","000000000000000101","111111111111110110","000000000000000000","111111111111101111","000000000000010100","000000000000000111","000000000000011000","000000000000100001","111111111111111001","111111111111101011","000000000000000000","111111111111110011","111111111111110101","000000000000000010","000000000000001011","000000000000001111","111111111111110011","111111111111110101","000000000000010011","111111111111011100","111111111111111100","111111111111111111","000000000000001100","111111111111101001","111111111111111110","111111111111011000","111111111111111010","000000000000001000","111111111111101110","000000000000000000","111111111111101101","111111111111111000","111111111111110000","000000000000000000","000000000000011011","000000000000011101","000000000000011100","111111111111101111","000000000000000010","000000000000000000","000000000000100001","111111111111100010","111111111111111101","000000000000000001","111111111111110100","000000000000010111","111111111111111110","000000000000000111","111111111111111111","111111111111101011","000000000000000110","111111111111101110","000000000000010010","000000000000000010","000000000000000001","000000000000001010","111111111111110001","000000000000001100","111111111111110110","000000000000001110","000000000000100001","111111111111100010","111111111111110001","000000000000010011","000000000000000011","000000000000000011","111111111111100110","111111111111111000","000000000000000001","000000000000000101","111111111111111001","111111111111101010","111111111111111010","000000000000001000","111111111111101001","111111111111111101","111111111111101111","000000000000001000","111111111111100010","111111111111101100","000000000000001101","000000000000100100","111111111111101101","000000000000011101","000000000000010011","000000000000000011","000000000000001010","111111111111011111","000000000000001000","000000000000010001","000000000000001110","000000000000100101","000000000000000000","000000000000010100","000000000000010011","000000000000000000","111111111111101110","000000000000000011","111111111111111100","111111111111101001","000000000000100001","111111111111110000","111111111111011111","111111111111100000","000000000000000101","000000000000010000","000000000000001101","111111111111011101","000000000000000000","000000000000000100","111111111111110111","111111111111111010","000000000000001101","111111111111110110","000000000000000000","000000000000000010","000000000000000100","000000000000000001","000000000000001010","000000000000000000","000000000000000110"),
("000000000000000011","000000000000000000","000000000000000011","111111111111110010","000000000000001000","111111111111110011","111111111111111110","000000000000010010","000000000000010001","111111111111110100","000000000000000000","000000000000001011","000000000000001010","000000000000000000","000000000000000000","111111111111111110","111111111111111100","111111111111101111","000000000000001111","111111111111110010","111111111111110001","000000000000000010","000000000000010100","000000000000001001","111111111111101101","000000000000000010","000000000000001001","000000000000001011","000000000000010001","000000000000001000","111111111111111100","000000000000001011","000000000000000000","111111111111111011","111111111111101111","111111111111110011","111111111111101100","000000000000001010","111111111111110011","111111111111101101","111111111111110000","111111111111111100","111111111111101110","000000000000000101","111111111111110001","000000000000010010","111111111111111010","111111111111110111","000000000000001010","111111111111101100","000000000000000000","000000000000000011","000000000000010000","111111111111110000","000000000000000010","000000000000010100","000000000000000011","111111111111111011","111111111111111100","111111111111110101","111111111111111010","111111111111111101","111111111111101101","111111111111111110","000000000000000100","000000000000001001","000000000000000011","000000000000010010","000000000000000100","111111111111110100","000000000000010010","111111111111111111","111111111111111000","000000000000010011","111111111111110000","000000000000000000","111111111111111110","000000000000000101","111111111111110100","000000000000001011","111111111111111101","000000000000000000","000000000000010011","111111111111110000","111111111111101101","000000000000000011","111111111111110001","111111111111110100","000000000000000000","000000000000000011","111111111111110010","111111111111111100","000000000000010011","000000000000001111","000000000000000011","000000000000000110","000000000000000110","000000000000000001","000000000000000010","111111111111101110","000000000000000000","111111111111110110","111111111111111010","111111111111111101","000000000000000001","000000000000001010","111111111111110000","000000000000000111","000000000000001101","111111111111110111","111111111111101101","111111111111110010","000000000000000001","000000000000001101","000000000000000101","111111111111111101","000000000000001000","000000000000000000","000000000000000001","111111111111110000","111111111111111011","111111111111110110","000000000000001101","000000000000010001","000000000000001010","111111111111101101","000000000000010000","111111111111101101"),
("000000000000001111","111111111111111101","111111111111110110","000000000000001100","000000000000000000","111111111111111110","000000000000010000","000000000000010100","111111111111110111","000000000000001111","111111111111101111","000000000000000100","111111111111111000","111111111111110010","000000000000000001","000000000000001001","000000000000010011","111111111111111111","000000000000000110","000000000000000011","111111111111110001","000000000000001011","111111111111110101","000000000000000110","111111111111101100","000000000000010001","111111111111110111","111111111111111001","000000000000001001","111111111111101101","111111111111110011","111111111111110110","111111111111110110","111111111111110101","000000000000000101","000000000000010000","000000000000010001","111111111111111111","111111111111111100","000000000000001011","000000000000001110","111111111111110100","111111111111111010","111111111111111000","000000000000010000","000000000000010011","000000000000000001","000000000000000100","000000000000010011","000000000000001000","000000000000001001","000000000000010000","111111111111110100","000000000000000000","000000000000001111","111111111111101111","000000000000000111","111111111111111010","000000000000001111","000000000000010001","111111111111111111","111111111111110111","111111111111110001","111111111111111010","000000000000001100","111111111111111000","000000000000000000","111111111111110100","000000000000010011","000000000000000100","111111111111110110","000000000000001111","000000000000000000","111111111111101111","111111111111110001","111111111111110011","000000000000000000","000000000000010011","111111111111110000","000000000000000110","000000000000000100","000000000000000000","000000000000000101","111111111111110011","111111111111101111","111111111111111100","000000000000000100","111111111111110011","000000000000001100","000000000000010100","000000000000001011","000000000000001000","000000000000001001","000000000000001101","000000000000010001","000000000000000101","111111111111111001","111111111111110000","000000000000000101","111111111111111110","000000000000000001","111111111111110101","000000000000000101","111111111111111011","000000000000001101","111111111111110010","111111111111110100","000000000000010001","000000000000001101","111111111111110110","000000000000000000","000000000000000110","000000000000010010","000000000000000011","000000000000000011","000000000000000011","111111111111111011","000000000000000111","000000000000001110","000000000000000101","000000000000000100","000000000000010100","111111111111110101","000000000000010001","111111111111101101","111111111111111101","000000000000000011","000000000000010010"),
("000000000000000010","111111111111110111","000000000000001000","111111111111111010","111111111111101111","000000000000001110","000000000000001101","111111111111111001","111111111111111100","000000000000000011","000000000000001101","000000000000010001","000000000000001111","111111111111111001","111111111111110000","000000000000000000","111111111111110101","000000000000000001","111111111111111110","111111111111110110","000000000000000111","111111111111110010","111111111111101101","111111111111111111","000000000000000001","111111111111110111","000000000000001101","111111111111101101","111111111111111011","111111111111111001","111111111111111101","000000000000010100","111111111111110001","111111111111110101","111111111111111010","111111111111101110","000000000000001001","111111111111110101","000000000000001101","111111111111111000","111111111111111110","111111111111111110","111111111111101101","000000000000010001","000000000000001011","000000000000010001","111111111111110111","111111111111111010","111111111111111101","000000000000000000","111111111111101100","000000000000001111","000000000000000000","000000000000000011","000000000000010011","000000000000000000","000000000000001100","000000000000010010","000000000000010001","000000000000000100","000000000000000000","000000000000001000","000000000000000111","000000000000000111","111111111111110001","000000000000000001","111111111111101100","000000000000001110","111111111111110100","000000000000000011","000000000000001011","000000000000010001","111111111111101101","000000000000001111","111111111111110001","111111111111110101","111111111111110011","111111111111111010","111111111111111001","000000000000001100","111111111111101111","111111111111111101","111111111111110111","000000000000000010","000000000000000001","111111111111101110","000000000000001100","000000000000001111","111111111111110111","000000000000010010","111111111111110001","111111111111101111","000000000000010001","000000000000010000","111111111111101101","111111111111111111","111111111111110000","111111111111110001","111111111111111001","000000000000010100","000000000000001011","000000000000000100","000000000000010010","000000000000000111","000000000000001001","111111111111101100","000000000000000000","111111111111111110","111111111111111111","000000000000001100","000000000000010010","111111111111110010","111111111111101100","000000000000010001","000000000000000111","111111111111110010","000000000000001101","111111111111110111","000000000000010001","000000000000010001","111111111111101110","111111111111111011","111111111111101101","000000000000001101","000000000000010010","000000000000000010","000000000000001101","111111111111110101"),
("111111111111110100","000000000000000100","000000000000000100","000000000000010010","111111111111101101","000000000000001111","000000000000010010","111111111111101110","000000000000000000","000000000000001111","000000000000000111","111111111111111010","000000000000010011","111111111111111000","111111111111111100","111111111111110100","000000000000010011","000000000000001101","000000000000001101","000000000000000101","111111111111110100","000000000000000010","000000000000000110","000000000000000100","000000000000000100","000000000000000010","000000000000000101","000000000000001101","000000000000000100","000000000000000100","111111111111111010","000000000000000100","111111111111110000","000000000000000000","000000000000010011","111111111111101101","000000000000000101","111111111111111001","000000000000001011","000000000000000010","111111111111111001","000000000000000010","111111111111110101","111111111111110100","111111111111101110","000000000000010000","111111111111111010","000000000000000110","000000000000001111","111111111111110100","000000000000001001","111111111111111110","111111111111110100","000000000000010010","111111111111111001","000000000000000100","000000000000001001","111111111111111101","111111111111101110","111111111111101111","000000000000001010","000000000000010010","111111111111111101","000000000000001011","000000000000000100","000000000000000110","111111111111110111","111111111111111001","111111111111110000","111111111111110011","000000000000001101","000000000000000110","000000000000000000","000000000000001110","111111111111111110","000000000000000100","111111111111110100","000000000000000100","111111111111111011","111111111111110011","000000000000000010","000000000000000000","111111111111110101","000000000000001101","000000000000000000","111111111111110101","000000000000010000","000000000000000100","111111111111110000","111111111111111010","111111111111111100","000000000000010100","000000000000001101","000000000000000000","000000000000010011","000000000000000011","000000000000000100","000000000000010000","111111111111110101","000000000000001010","111111111111111111","111111111111101111","111111111111111101","000000000000000010","000000000000000000","000000000000000100","111111111111110100","111111111111111001","000000000000010100","000000000000000111","000000000000000111","111111111111111110","000000000000000100","111111111111101110","111111111111111101","111111111111110100","111111111111110101","000000000000000010","111111111111111110","111111111111110000","111111111111110010","111111111111111000","000000000000000110","000000000000010100","111111111111110000","111111111111101110","000000000000001110","000000000000000101"),
("111111111111111011","111111111111111101","000000000000000001","111111111111110001","111111111111101111","000000000000010000","111111111111110000","000000000000001001","111111111111111100","000000000000001011","111111111111110001","111111111111111111","111111111111110000","000000000000000001","000000000000001101","111111111111111000","000000000000001011","111111111111110001","111111111111111010","000000000000001010","111111111111111111","000000000000010000","000000000000001010","111111111111110010","000000000000000011","111111111111110111","000000000000010000","111111111111110111","111111111111101101","000000000000010100","111111111111110101","000000000000001001","111111111111110001","111111111111101110","000000000000000100","000000000000000000","000000000000000010","111111111111101110","000000000000000110","111111111111111010","000000000000001110","111111111111101110","000000000000000000","111111111111101110","000000000000001001","111111111111110011","111111111111101101","000000000000001010","111111111111111011","000000000000000101","111111111111110010","000000000000000011","111111111111111101","111111111111111000","000000000000000101","111111111111111101","111111111111110100","000000000000001101","000000000000001111","111111111111110110","000000000000001010","000000000000000010","111111111111111100","111111111111101100","111111111111110001","111111111111111001","111111111111110101","000000000000001101","000000000000001100","000000000000000000","111111111111101101","000000000000001001","000000000000001110","000000000000010100","111111111111110010","111111111111111000","000000000000001110","111111111111110001","111111111111110110","111111111111111000","000000000000000010","000000000000000000","000000000000000110","000000000000010010","000000000000000000","000000000000001100","000000000000001010","111111111111111001","111111111111111100","000000000000000001","000000000000000001","000000000000010011","000000000000000000","111111111111110111","111111111111110100","000000000000000001","111111111111101101","000000000000010010","111111111111111101","000000000000010011","111111111111110001","111111111111111001","111111111111110101","111111111111110100","111111111111101100","000000000000010000","000000000000000111","111111111111111110","111111111111111001","000000000000000001","111111111111110101","111111111111110010","000000000000001100","000000000000001010","000000000000000101","111111111111110101","111111111111110100","000000000000010100","111111111111101111","111111111111111100","000000000000000110","000000000000001000","111111111111110001","111111111111110001","000000000000000000","000000000000000001","000000000000010010","111111111111101110"),
("000000000000000101","111111111111111000","111111111111110010","111111111111110110","111111111111111001","000000000000001101","111111111111110011","111111111111111100","000000000000010010","000000000000001001","000000000000000111","111111111111110110","000000000000001011","000000000000000001","000000000000010100","111111111111110100","111111111111111001","000000000000001001","111111111111111010","111111111111110100","000000000000010010","000000000000001111","000000000000000000","000000000000000101","111111111111110011","000000000000000111","000000000000000000","111111111111110111","111111111111110010","111111111111111100","111111111111110001","111111111111110111","111111111111101110","000000000000000100","000000000000000101","000000000000001010","111111111111111001","111111111111111101","111111111111111110","111111111111111011","000000000000010000","000000000000000111","111111111111111001","111111111111101101","111111111111111110","111111111111101100","000000000000000000","000000000000000000","000000000000010001","000000000000001101","111111111111101101","111111111111110111","111111111111110000","111111111111111011","111111111111110000","111111111111101110","000000000000001001","111111111111101111","000000000000000111","111111111111101101","111111111111110001","111111111111110100","000000000000010000","000000000000001001","000000000000000000","111111111111110011","111111111111111101","000000000000000010","000000000000001100","000000000000001101","111111111111110001","000000000000000100","000000000000010011","111111111111111100","000000000000001001","111111111111111000","000000000000000011","111111111111110001","000000000000000011","111111111111101111","111111111111110000","111111111111110110","111111111111110000","111111111111111000","111111111111110110","111111111111111110","000000000000000111","000000000000001000","000000000000000110","111111111111111101","000000000000010011","000000000000001011","111111111111110011","000000000000001001","000000000000000100","000000000000000110","000000000000001111","000000000000010000","111111111111110011","111111111111111001","000000000000010010","000000000000001101","111111111111110111","000000000000000000","000000000000000000","111111111111110101","000000000000000100","111111111111110010","111111111111110001","000000000000000010","111111111111110000","111111111111110000","000000000000000010","000000000000000000","111111111111110100","111111111111111010","111111111111110110","000000000000010001","000000000000001010","111111111111110010","000000000000001000","111111111111111111","000000000000000101","111111111111110010","000000000000001010","000000000000000111","000000000000001101","000000000000001100"),
("111111111111110001","000000000000001111","111111111111111010","000000000000000000","111111111111110101","111111111111101110","000000000000010100","000000000000010010","000000000000001110","000000000000000101","000000000000001001","111111111111110100","111111111111111011","111111111111110111","111111111111111110","000000000000010100","111111111111101101","111111111111110100","111111111111110111","000000000000000000","000000000000010001","000000000000000001","000000000000000010","000000000000000110","000000000000000001","000000000000001101","000000000000001011","000000000000000111","000000000000000001","000000000000000010","111111111111111000","000000000000001001","000000000000000011","111111111111110111","111111111111110101","000000000000001000","111111111111101101","111111111111101101","000000000000001000","000000000000001001","111111111111101110","000000000000010001","000000000000001011","111111111111110000","111111111111110011","000000000000000000","000000000000000111","000000000000010100","111111111111110111","000000000000000000","000000000000001101","000000000000001110","000000000000010010","000000000000000000","000000000000000111","111111111111110010","000000000000010000","111111111111111001","000000000000001111","000000000000010010","000000000000001100","111111111111111000","000000000000010010","111111111111110001","111111111111111000","111111111111111011","111111111111111111","111111111111110001","111111111111111100","000000000000000001","000000000000010010","111111111111110101","000000000000001001","111111111111101100","000000000000010000","111111111111111111","111111111111110100","000000000000001101","111111111111110100","111111111111101111","111111111111111011","111111111111101111","111111111111111101","111111111111111000","000000000000001110","000000000000000000","000000000000000001","000000000000001011","000000000000001001","000000000000000000","000000000000001001","000000000000000101","111111111111101111","000000000000010100","000000000000000111","111111111111101111","111111111111110110","000000000000001111","000000000000010001","000000000000001001","000000000000000101","000000000000000000","000000000000010011","000000000000010001","000000000000010000","111111111111110110","000000000000001100","000000000000000010","111111111111110111","111111111111110110","000000000000010000","111111111111111011","111111111111111011","111111111111111101","000000000000000010","000000000000000011","111111111111101111","000000000000000100","111111111111111011","111111111111111110","000000000000001110","111111111111110100","000000000000010101","000000000000001101","000000000000000011","000000000000000111","000000000000000100","000000000000000011"),
("111111111111111000","000000000000000101","111111111111110001","000000000000011010","000000000000010010","000000000000000000","000000000000000100","000000000000001110","111111111111110110","000000000000000001","000000000000001110","000000000000010110","000000000000001110","000000000000000001","111111111111111001","000000000000001110","111111111111111011","111111111111110100","000000000000001000","111111111111111000","000000000000001000","000000000000001010","000000000000010110","000000000000011011","111111111111111110","111111111111100110","111111111111100101","000000000000010001","111111111111111101","000000000000001100","111111111111101100","111111111111111011","000000000000000000","000000000000001001","111111111111111110","111111111111101100","111111111111100110","000000000000000101","111111111111110100","111111111111100100","000000000000001011","000000000000010000","111111111111101110","111111111111111111","111111111111110111","000000000000001110","111111111111111100","111111111111101111","111111111111110001","111111111111100111","000000000000011000","000000000000000111","000000000000001011","111111111111111001","000000000000001000","111111111111100101","111111111111110000","000000000000010010","000000000000010111","000000000000010010","000000000000011101","111111111111110111","111111111111111111","111111111111101100","000000000000000000","000000000000001001","000000000000000110","000000000000101000","000000000000001000","111111111111111000","111111111111110001","000000000000000100","000000000000001111","111111111111101101","111111111111110011","000000000000001111","111111111111011110","000000000000000101","111111111111111101","111111111111101000","111111111111111101","111111111111111001","111111111111110010","111111111111101100","000000000000001111","111111111111110011","000000000000000111","111111111111110100","000000000000000011","000000000000010010","111111111111100101","000000000000011010","000000000000001001","000000000000000110","000000000000010000","111111111111110101","000000000000001001","111111111111110010","111111111111101010","111111111111011111","000000000000001010","111111111111101110","000000000000011011","000000000000011011","111111111111110110","000000000000100010","111111111111100001","111111111111101010","111111111111101011","000000000000000100","111111111111110001","000000000000010001","111111111111101001","000000000000001010","111111111111111001","000000000000100100","000000000000101001","111111111111110001","000000000000001000","000000000000000100","000000000000001110","000000000000010101","111111111111110101","000000000000000101","000000000000011110","111111111111110111","111111111111110111","111111111111110101"),
("111111111111111101","000000000000100010","000000000000000110","111111111111110100","111111111111101111","000000000000000001","000000000000000010","000000000000001011","000000000000001010","000000000000010011","000000000000001011","000000000000000100","000000000000000110","111111111111110100","111111111111100000","000000000000000000","000000000000000010","111111111111110110","000000000000001100","000000000000001111","000000000000001110","000000000000010011","111111111111111011","111111111111101101","000000000000010011","111111111111110101","111111111111100000","000000000000001110","111111111111110001","111111111111111000","111111111111100110","111111111111111100","000000000000010110","000000000000000001","111111111111101001","111111111111111101","000000000000000000","111111111111111100","111111111111101110","111111111111111010","111111111111111100","000000000000011111","000000000000011010","000000000000001100","111111111111111111","111111111111110001","111111111111111001","111111111111100111","111111111111011110","111111111111111110","000000000000000010","000000000000001011","000000000000100001","111111111111110010","111111111111111000","111111111111101001","000000000000001010","111111111111111111","000000000000011001","111111111111110000","000000000000011011","111111111111101110","111111111111110101","111111111111101011","000000000000000101","000000000000010010","111111111111111100","000000000000000011","111111111111111010","000000000000000101","000000000000010111","000000000000010010","000000000000011000","111111111111101101","000000000000000110","111111111111110100","111111111111101101","000000000000001101","111111111111101110","111111111111110110","000000000000001010","000000000000000110","000000000000000010","000000000000001000","000000000000000100","000000000000000001","000000000000000111","111111111111110111","111111111111111010","000000000000001011","000000000000001111","000000000000000101","000000000000001011","000000000000000011","111111111111111100","111111111111110100","111111111111111001","111111111111110111","000000000000000010","111111111111100001","111111111111110011","111111111111101000","111111111111110111","000000000000001101","111111111111110110","000000000000100010","111111111111100100","000000000000001011","000000000000000010","000000000000000011","000000000000001011","000000000000000011","111111111111110100","111111111111101010","111111111111100011","000000000000010010","000000000000001101","000000000000010010","111111111111101101","111111111111111100","000000000000001110","000000000000000111","111111111111110110","000000000000010011","000000000000000100","111111111111111101","111111111111110001","111111111111111001"),
("000000000000000100","000000000000000011","000000000000001000","000000000000001011","111111111111111100","000000000000001110","000000000000010001","000000000000000111","000000000000000001","111111111111110000","000000000000000000","111111111111111010","111111111111111100","000000000000001110","000000000000011010","000000000000001100","000000000000001010","111111111111110001","000000000000001000","000000000000000100","111111111111101100","111111111111110110","000000000000001000","000000000000001100","111111111111110001","000000000000010111","000000000000001000","111111111111111000","000000000000001111","111111111111110101","000000000000010100","000000000000001000","111111111111110111","000000000000001101","111111111111110010","111111111111110011","000000000000001101","000000000000000110","000000000000000101","111111111111101111","000000000000001010","111111111111110101","000000000000100111","000000000000100111","111111111111110011","111111111111101110","000000000000011000","000000000000011001","111111111111100011","000000000000000000","000000000000000111","000000000000001100","111111111111111111","000000000000000100","111111111111100010","111111111111111111","111111111111111101","000000000000001110","000000000000000100","000000000000000101","111111111111111111","000000000000001110","111111111111110110","111111111111111101","111111111111111101","111111111111110011","111111111111111010","000000000000001001","000000000000000101","000000000000000000","000000000000001000","111111111111111101","111111111111111111","111111111111111110","000000000000011010","000000000000010001","111111111111110111","111111111111101100","111111111111101110","000000000000001010","000000000000010101","000000000000010010","111111111111101111","111111111111111101","000000000000001000","000000000000010010","000000000000010001","000000000000001111","000000000000010000","111111111111111010","111111111111111001","111111111111110100","111111111111110110","000000000000000010","111111111111110111","111111111111111011","111111111111101101","000000000000011010","000000000000010010","111111111111111111","000000000000001010","111111111111111110","000000000000001101","000000000000010001","111111111111111010","000000000000000100","111111111111110111","111111111111110110","111111111111101010","000000000000010101","111111111111101100","111111111111110000","000000000000000001","111111111111101101","111111111111111011","000000000000010010","000000000000000111","111111111111110100","000000000000001000","111111111111100011","111111111111110011","000000000000000000","111111111111111010","111111111111111001","000000000000001011","111111111111101111","000000000000011011","111111111111101001"),
("000000000000001100","000000000000011111","111111111111011110","111111111111110010","000000000000000001","000000000000000101","000000000000001110","111111111111100101","000000000000000101","000000000000001000","111111111111111111","000000000000100000","000000000000010011","000000000000000101","000000000000011100","000000000000000101","111111111111111000","000000000000000000","000000000000001111","000000000000000000","000000000000000001","111111111111011100","111111111111100000","000000000000010000","111111111111101110","000000000000010101","111111111111111100","111111111111101111","000000000000001011","000000000000001010","000000000000001000","000000000000010110","111111111111101111","111111111111111010","000000000000001110","111111111111100011","000000000000010000","111111111111111110","111111111111100001","111111111111110110","000000000000000000","000000000000001011","000000000000011100","000000000000001000","111111111111111010","000000000000000010","000000000000101101","000000000000001100","111111111111100111","000000000000011100","111111111111110010","111111111111101000","111111111111110000","111111111111011110","111111111111110010","111111111111110010","000000000000000100","111111111111110001","111111111111100000","111111111111110000","111111111111111010","111111111111101010","111111111111110101","111111111111100110","111111111111101101","111111111111110011","000000000000001010","000000000000011011","111111111111011110","111111111111110001","000000000000011101","111111111111110010","000000000000011001","111111111111100111","000000000000010110","000000000000000110","000000000000000100","000000000000001010","111111111111110011","111111111111110111","000000000000000111","111111111111101000","111111111111111100","111111111111111111","000000000000000000","111111111111111011","111111111111011101","000000000000011010","111111111111111111","000000000000000110","000000000000010111","111111111111110010","000000000000011111","000000000000000011","111111111111011100","000000000000000000","000000000000001100","000000000000011100","000000000000001110","111111111111111011","000000000000011110","000000000000010000","000000000000010111","111111111111111011","111111111111110101","000000000000011001","111111111111100010","000000000000010010","111111111111100010","111111111111101101","111111111111011010","111111111111110011","000000000000100000","111111111111110110","111111111111110100","000000000000000111","000000000000000010","000000000000001000","111111111111110111","111111111111110001","000000000000000000","111111111111111111","000000000000001100","000000000000110110","000000000000001111","000000000000010010","000000000000001111","000000000000000000"),
("000000000000001010","000000000000001110","111111111111011100","000000000000001110","111111111111111001","111111111111110101","000000000000011101","111111111111101100","111111111111100010","000000000000100101","000000000000000000","000000000000100010","111111111111111010","000000000000000100","000000000000010001","000000000000001110","111111111111101011","111111111111111011","000000000000001000","111111111111111011","000000000000001010","000000000000011010","111111111111100101","000000000000010111","111111111111111011","000000000000001111","111111111111110010","111111111111110001","000000000000001100","111111111111111010","111111111111111100","000000000000011010","111111111111110010","111111111111111010","111111111111111010","111111111111101101","111111111111110001","111111111111111011","111111111111111000","111111111111101100","111111111111110100","000000000000000111","000000000000000110","000000000000001111","111111111111010110","000000000000000001","000000000000100011","000000000000000000","111111111111101101","111111111111111100","111111111111101100","111111111111011100","000000000000010111","111111111111011111","111111111111101100","111111111111100101","000000000000000011","111111111111101101","111111111111111111","111111111111110100","000000000000001001","000000000000001001","111111111111101100","111111111111101001","111111111111101110","111111111111101100","000000000000001010","000000000000001101","111111111111011011","111111111111101010","000000000000001100","111111111111101100","000000000000001010","111111111111100001","000000000000100110","000000000000001101","111111111111100000","000000000000001001","111111111111011110","111111111111110111","111111111111111110","111111111111100000","000000000000000100","111111111111111101","111111111111110000","000000000000000010","111111111111101000","000000000000000100","000000000000011010","111111111111111101","000000000000001000","000000000000001011","000000000000100011","000000000000010100","111111111111110000","111111111111111011","111111111111101011","000000000000010100","000000000000000001","111111111111101001","000000000000010010","000000000000011000","111111111111111111","000000000000000000","000000000000010010","000000000000011101","111111111111100111","000000000000011000","111111111111110010","111111111111110001","111111111111011101","111111111111101110","000000000000000110","111111111111110001","111111111111101111","000000000000010111","000000000000010011","111111111111100100","111111111111110111","000000000000000011","111111111111111001","000000000000010101","000000000000100001","000000000000011100","000000000000011111","000000000000001001","000000000000010011","111111111111100000"),
("111111111111111010","000000000000001100","111111111111111000","000000000000000000","000000000000010110","000000000000100110","000000000000010000","000000000000000101","000000000000000011","000000000000000001","000000000000010100","000000000000000010","111111111111111101","000000000000001011","000000000000010001","000000000000100010","111111111111110010","111111111111110000","000000000000000001","111111111111100111","111111111111111010","000000000000000110","111111111111010001","111111111111101100","000000000000000011","000000000000101110","111111111111111010","000000000000011011","000000000000101001","000000000000010110","111111111111110110","000000000000101000","111111111111110001","000000000000001000","000000000000110010","111111111111100000","000000000000011010","000000000000000011","111111111111101010","111111111111101010","111111111111111011","111111111111110110","000000000000101011","000000000000100111","111111111111111001","111111111111101001","000000000000011000","000000000000101000","111111111111011111","000000000000001101","111111111111101110","111111111111101010","000000000000010000","111111111111011010","000000000000000101","111111111111010011","111111111111110011","111111111111111100","111111111111101100","111111111111110000","000000000000000101","000000000000001100","000000000000000110","111111111111101001","111111111111111010","111111111111110111","000000000000010110","000000000000100101","000000000000000000","111111111111100010","000000000000001100","000000000000001000","000000000000010000","111111111111011010","000000000000000010","000000000000010010","111111111111110101","000000000000000000","000000000000000000","000000000000000010","000000000000001000","000000000000000001","000000000000000101","111111111111101101","111111111111011011","000000000000000100","111111111111101100","000000000000010101","111111111111111001","111111111111101010","000000000000000100","111111111111101111","000000000000110000","000000000000011001","111111111111101001","111111111111111110","000000000000000010","000000000000100111","111111111111110001","111111111111111100","000000000000001100","000000000000010011","000000000000011000","000000000000000010","000000000000000010","000000000000010100","111111111111011111","000000000000001110","000000000000000000","111111111111111111","111111111111100101","111111111111110111","000000000000010100","111111111111011010","111111111111010000","000000000000010011","000000000000011000","111111111111100101","111111111111110011","000000000000000000","000000000000001000","000000000000000001","000000000000001100","000000000000010001","000000000000010111","000000000000000000","000000000000011110","111111111111011111"),
("111111111111111011","111111111111111111","111111111111001111","000000000000010000","000000000000101001","000000000000100110","000000000000010000","000000000000001010","000000000000000101","111111111111111010","000000000000010100","111111111111111011","111111111111101110","000000000000000000","000000000000101100","000000000000101010","000000000000000101","111111111111110101","111111111111111111","000000000000001110","111111111111101101","111111111111110000","111111111111110011","000000000000000010","111111111111101011","000000000001000010","111111111111010011","000000000000001111","000000000000011000","111111111111110011","000000000000011111","000000000000010000","111111111111111111","111111111111110110","000000000000111100","111111111111110100","000000000000001000","000000000000000011","111111111111101110","111111111111011011","000000000000000011","111111111111101010","000000000000101001","000000000000110110","111111111111111111","111111111111101010","000000000000001000","000000000000101001","111111111111000110","000000000000011110","000000000000000001","111111111111111011","111111111111101111","111111111111110110","111111111111111011","111111111111101000","111111111111110011","111111111111011101","111111111111010101","111111111111111010","111111111111100110","000000000000011100","111111111111111000","111111111111100110","000000000000000000","111111111111100101","111111111111110000","000000000000000000","000000000000000110","111111111111111110","000000000000110100","000000000000011001","000000000000001010","000000000000001011","000000000000000100","000000000000101000","000000000000001001","000000000000001001","000000000000010010","111111111111110011","111111111111100100","000000000000000101","000000000000111100","111111111111111100","111111111111101111","111111111111100101","111111111111101111","000000000000001101","111111111111111111","000000000000000111","111111111111101011","111111111111101011","000000000000000111","000000000000000110","111111111111100011","000000000000010010","111111111111110111","000000000000010011","111111111111010000","000000000000000101","000000000000010111","111111111111111101","000000000000000000","111111111111111011","111111111111011111","000000000000101111","111111111111100101","000000000000000101","111111111111110000","111111111111100010","111111111111101011","111111111111110010","000000000000010010","111111111111101111","111111111111100110","000000000000010111","000000000000000110","000000000000001111","111111111111100101","000000000000100011","000000000000101101","000000000000001011","000000000000011011","000000000000100100","000000000000110001","111111111111110000","000000000000100011","111111111111111001"),
("000000000000000000","000000000000010011","111111111111011110","000000000000000001","000000000000001011","000000000000010011","000000000000110001","000000000000000000","000000000000010101","000000000000100001","000000000000010000","111111111111111010","000000000000001010","111111111111110001","000000000000011001","000000000000101010","000000000000001110","111111111111111111","000000000000011111","111111111111110101","111111111111100010","111111111111001100","111111111111101101","111111111111101011","111111111111111000","000000000000111101","111111111111010111","000000000000000001","000000000000100000","111111111111110110","000000000000000001","000000000000010010","000000000000010010","111111111111101111","000000000000100000","111111111111110000","000000000000010110","000000000000000111","111111111111001001","111111111111101110","111111111111111101","111111111111101001","000000000000100110","000000000000101101","111111111111111000","111111111111001010","000000000000100110","000000000000011111","111111111110111100","000000000000000010","111111111111110010","111111111111111111","111111111111111101","111111111111111111","000000000000000101","000000000000000000","111111111111010110","111111111111100011","111111111111010110","111111111111110010","111111111111110111","000000000000001110","000000000000000100","111111111111101110","111111111111011010","111111111111001000","111111111111110100","000000000000000110","000000000000001010","111111111111111101","000000000000100110","000000000000000110","111111111111111111","000000000000010110","000000000000000100","000000000000100101","000000000000000010","000000000000000100","111111111111100111","111111111111110101","111111111111010011","000000000000000100","000000000000100011","111111111111011010","111111111111110010","111111111111110111","111111111111101001","111111111111111010","111111111111111000","000000000000001000","111111111111111111","111111111111101100","000000000000011100","000000000000011100","111111111111011000","111111111111111101","000000000000011111","000000000000100011","111111111111100010","111111111111011101","000000000000111011","000000000000010110","000000000000001111","000000000000001111","111111111111100011","000000000000011011","111111111111010000","000000000000101001","111111111111110110","111111111111110101","111111111111101110","111111111111100100","000000000000000110","111111111111101110","111111111111010011","000000000000011111","000000000000010101","111111111111110101","111111111111010001","000000000000101100","000000000000011100","000000000000001000","000000000000111001","000000000000011101","000000000000010010","000000000000000011","000000000000111001","111111111111101000"),
("000000000000000001","000000000000101101","111111111111011010","000000000000001011","000000000000000000","000000000000011011","000000000000111000","111111111111111001","000000000000010101","000000000000110000","000000000000001011","000000000000011111","000000000000010010","000000000000000111","000000000000100011","000000000000011001","000000000000010111","111111111111110111","000000000000001100","000000000000010110","111111111111010000","111111111111100000","111111111111000110","111111111111100100","111111111111011111","000000000000110011","111111111111110010","000000000000100110","000000000000001000","000000000000000111","000000000000001000","000000000000000001","000000000000010010","000000000000001100","111111111111111000","111111111111110110","000000000000010110","111111111111111000","111111111111100001","111111111111101000","111111111111010000","111111111111111010","000000000001010100","000000000001001111","000000000000000010","111111111111011110","000000000000101011","000000000000001111","111111111111000110","111111111111111010","000000000000010101","000000000000000000","111111111111101100","111111111111101001","000000000000000000","111111111111111100","111111111111010111","111111111111110010","111111111111100000","111111111111111100","000000000000000011","000000000000010110","111111111111110000","111111111111100110","111111111111110100","111111111111001010","111111111111110001","000000000000011100","000000000000000011","111111111111110011","000000000001001110","000000000000010100","111111111111100000","000000000000001001","000000000000010111","000000000000101011","111111111111101010","000000000000001010","000000000000000110","000000000000000011","111111111111100001","111111111111111111","000000000000001110","111111111111011100","111111111111110110","111111111111100011","111111111111110000","000000000000010111","000000000000011001","111111111111111110","000000000000000011","000000000000001100","000000000000011001","000000000000001011","111111111110111011","111111111111100111","000000000000000000","000000000000110101","111111111111100011","111111111111101010","000000000000001010","000000000000000100","111111111111110100","000000000000000001","000000000000000100","000000000000111101","111111111111101100","000000000000110000","111111111111011101","111111111111111101","111111111111100011","111111111111110010","000000000000001101","111111111111111000","111111111110101101","000000000000101011","000000000000110101","111111111111100011","111111111111111001","000000000000001101","000000000000000110","111111111111110000","000000000000111010","111111111111110101","000000000000101011","111111111111111100","000000000000011101","111111111111100010"),
("111111111111111001","000000000000011111","111111111111101100","000000000000000110","111111111111010010","000000000000010011","000000000000100111","000000000000000111","111111111111110101","000000000000000111","000000000000000000","000000000000000000","000000000000010101","111111111111101110","000000000000101101","000000000000110010","000000000000011101","000000000000010001","000000000000010110","000000000000000101","111111111111101001","111111111111101000","111111111111010010","111111111111110110","111111111111011011","000000000000100001","111111111111010101","000000000000010011","000000000000001100","000000000000000101","000000000000010001","000000000000011110","000000000000000010","111111111111110110","000000000000011001","111111111111111101","000000000000000010","000000000000000101","111111111111110101","111111111111110001","111111111111110010","111111111111100111","000000000000100001","000000000000100011","111111111111011001","111111111111011100","000000000000011101","000000000000100001","111111111111100110","111111111111111001","111111111111110110","111111111111110111","111111111111111001","111111111111100110","000000000000001111","111111111111011111","111111111111110011","000000000000001110","111111111111100100","111111111111110100","111111111111111110","000000000000100010","000000000000010101","111111111111011101","111111111111110010","111111111111010010","111111111111101110","000000000000011100","111111111111110000","111111111111100010","000000000000101010","000000000000100110","000000000000000000","000000000000000101","000000000000000100","000000000000011111","000000000000000100","000000000000011101","000000000000000000","111111111111110100","111111111111101000","000000000000010101","000000000000010010","111111111111010111","000000000000001001","000000000000001000","111111111111011100","000000000000101000","000000000000001011","111111111111111001","111111111111111110","000000000000010110","000000000000010110","000000000000011101","111111111111010010","111111111111011000","000000000000000000","000000000000001101","111111111111010011","111111111111100100","000000000000011011","000000000000001110","000000000000010100","111111111111111001","000000000000000001","000000000000101110","111111111111001111","000000000000010010","111111111111000111","111111111111110100","111111111110111110","111111111111011100","000000000000011110","000000000000000100","111111111110101010","000000000000010101","000000000000001100","111111111111110011","111111111111001101","000000000000001000","111111111111111110","111111111111111100","000000000000100111","000000000000010010","000000000000010001","000000000000011101","000000000000100011","111111111111010101"),
("111111111111101111","000000000000011111","111111111111100001","000000000000100000","111111111111010001","000000000000010100","111111111111111110","111111111111110110","111111111111110111","111111111111101011","000000000000001100","111111111111101010","111111111111110001","111111111111100000","000000000000100100","111111111111110111","000000000000111110","111111111111111000","111111111111110000","000000000000001001","000000000000011001","111111111111110001","000000000000000001","111111111111011101","111111111111010101","000000000000001100","111111111111011100","000000000000001100","000000000000101100","111111111111111011","111111111111110110","000000000000101100","111111111111100100","000000000000100000","000000000000010110","111111111111010001","111111111111110000","111111111111111101","000000000000000000","111111111111100011","000000000000001011","111111111111101101","000000000000101111","000000000000100101","111111111111011000","000000000000000000","000000000000000100","000000000001000111","111111111111001000","111111111111111011","111111111111101101","111111111111110000","111111111111101101","111111111111111100","000000000000010110","111111111111110100","111111111111110101","111111111111111101","111111111111001101","000000000000001110","111111111111100111","000000000000011011","000000000000100011","000000000000000000","111111111111111000","111111111111010111","111111111111100000","000000000000000001","111111111111101010","111111111111101010","000000000000110110","000000000000010001","111111111111001010","111111111111111101","000000000000011000","000000000000000000","111111111111100010","000000000000011001","111111111111110000","111111111111111101","111111111111100100","111111111111011100","000000000000001111","111111111111010010","000000000000011000","000000000000000100","111111111111111000","000000000000001011","111111111111111010","111111111111111110","000000000000101001","111111111111101001","111111111111111110","000000000000101110","111111111111001111","000000000000010000","111111111111110001","111111111111110100","111111111111100000","000000000000001010","111111111111111001","000000000000101010","111111111111101111","000000000000010101","111111111111111011","000000000000000101","111111111111000110","000000000000001001","111111111111010110","111111111111111101","111111111111100110","111111111111011110","111111111111110000","111111111111011000","111111111110111011","000000000000001110","111111111111110011","111111111111111011","111111111110111100","000000000000001001","000000000000000010","000000000000001010","000000000000100010","000000000000101101","000000000000000010","000000000000000011","111111111111111110","111111111111110001"),
("000000000000001011","000000000000001011","111111111111010010","000000000000001100","111111111111000010","000000000000100111","000000000000010110","111111111111101101","111111111111111101","111111111111100011","000000000000011000","111111111111101011","111111111111100110","111111111111010000","000000000000110000","000000000000001100","000000000000100010","111111111111110110","111111111111111101","000000000000001101","111111111111111100","000000000000000000","000000000000001100","111111111111101101","111111111111011110","000000000000101110","111111111111100001","111111111111111111","000000000000010100","111111111111101000","000000000000011101","000000000000011110","111111111111101010","111111111111111001","000000000000100011","111111111111010110","111111111111110101","111111111111110110","111111111111101110","000000000000000000","000000000000011001","000000000000000001","000000000000111011","000000000001010001","111111111111101010","111111111111101110","000000000000101100","000000000000100001","111111111111101000","111111111111111111","111111111111111011","111111111111110100","111111111111000010","111111111111101110","000000000000001000","000000000000000000","000000000000001001","111111111111110110","111111111111011010","111111111111111011","111111111111010111","000000000000100110","000000000000011100","000000000000001000","111111111111111000","111111111111000111","111111111111000000","111111111111111111","111111111111010010","111111111111110010","000000000000100010","000000000000000111","111111111111010001","111111111111101100","000000000000101001","000000000000000111","000000000000011110","000000000000000111","000000000000011000","111111111111110010","000000000000000000","111111111111100100","000000000000011110","111111111111000101","000000000000001011","000000000000000111","111111111111100110","000000000000100101","111111111111110110","111111111111111110","000000000000010011","111111111111101001","000000000000001010","000000000000010010","111111111111001000","000000000000111001","000000000000000001","111111111111101010","111111111111101101","111111111111101011","111111111111111111","000000000000101100","111111111111101111","000000000000000100","111111111111110110","000000000000010011","111111111111001001","000000000000110010","111111111111010100","111111111111110001","111111111111100100","111111111111110010","000000000000010101","111111111111101001","111111111111101100","000000000000010110","000000000000000011","111111111111111011","111111111111000101","111111111111101101","111111111111110100","000000000000001100","000000000000111010","000000000000010101","000000000000100111","000000000000010110","000000000000100100","111111111111101100"),
("111111111111111010","000000000000001110","111111111111010110","000000000000011000","111111111110100011","000000000000001010","000000000000000100","111111111111010101","000000000000000010","000000000000001011","000000000000001011","111111111111111101","000000000000000011","111111111111011110","000000000001000010","000000000000100000","000000000000100001","111111111111111011","111111111111101110","111111111111100100","000000000000001010","111111111111100000","111111111111101010","111111111111111001","111111111111010100","000000000000010100","111111111111111110","111111111111111000","000000000000101111","111111111111100011","000000000000100101","000000000000101010","111111111111010111","000000000000010111","000000000000011010","000000000000000010","111111111111100001","000000000000001011","111111111111010101","111111111111111100","000000000000100111","000000000000011001","000000000000001011","000000000001001000","111111111111000111","000000000000011111","000000000000010000","000000000000101010","111111111111011001","111111111111110000","000000000000000100","111111111111011101","111111111111101010","000000000000000000","000000000000000110","111111111111111100","000000000000010100","111111111111111001","111111111110110111","111111111111110000","111111111111101001","000000000000011111","000000000000010111","111111111111110000","000000000000000100","111111111111010010","111111111111001101","000000000000010100","111111111111110100","111111111111111000","000000000001000011","000000000000010000","111111111111000011","111111111111010001","000000000000110010","000000000000000001","000000000000000010","000000000000001111","000000000000010111","111111111111110001","000000000000000000","111111111111110111","000000000000001101","111111111111001000","000000000000000101","111111111111100100","111111111111100011","000000000000100111","111111111111111101","000000000000101000","000000000000010100","111111111111011100","111111111111101101","000000000000011111","111111111110101001","000000000000110101","111111111111011001","000000000000001111","000000000000010011","111111111111100100","111111111111110100","000000000000011110","000000000000000101","000000000000011000","000000000000001001","000000000000001110","111111111111001100","000000000000001100","111111111111011000","111111111111111101","111111111111100011","111111111111101011","000000000000001100","111111111111101001","111111111111100011","111111111111111000","000000000000000111","111111111111110001","111111111111000001","111111111111111001","000000000000000010","000000000000000100","000000000000110001","111111111111101001","000000000000010010","000000000000010101","111111111111111011","111111111111010001"),
("111111111111101101","000000000000001101","111111111111100101","000000000000001001","111111111111000001","111111111111111101","111111111111111110","111111111111100011","111111111111110001","000000000000011001","111111111111110000","000000000000010000","000000000000100000","111111111111000011","000000000000011011","000000000000011100","000000000000010011","000000000000011101","111111111111100111","111111111111101011","000000000000000011","111111111111100110","111111111111011101","111111111111110010","111111111111111000","000000000000010110","111111111111110111","111111111111110101","000000000000100011","000000000000011001","000000000000000101","000000000000101101","111111111111010110","000000000000101000","000000000000101000","111111111111111100","000000000000001010","000000000000011101","111111111111011011","111111111111111100","000000000000110101","000000000000101011","000000000000001010","000000000000000111","111111111111010110","000000000000011011","000000000000011010","000000000000010100","111111111111011010","111111111111101110","111111111111110001","111111111111100001","000000000000000111","000000000000010000","000000000000010011","111111111111110100","111111111111111011","111111111111100100","111111111111000001","111111111111110111","000000000000010100","000000000000010101","000000000000000110","111111111111011001","111111111111101100","111111111111001011","111111111111010100","000000000000010011","111111111111100111","111111111111111101","000000000000101110","000000000000010110","111111111111100100","111111111111011000","000000000000011111","111111111111101100","111111111111110110","111111111111110111","111111111111101000","111111111111100010","111111111111101010","111111111111010010","000000000000000110","111111111110111100","000000000000001100","111111111111011111","111111111111110110","000000000000100110","000000000000000101","111111111111110110","111111111111111110","111111111111100010","111111111111110111","000000000000101011","111111111111000100","000000000000101001","111111111111101000","111111111111111001","000000000000011111","111111111111110000","111111111111110111","111111111111111001","111111111111110101","000000000000010010","111111111111111011","111111111111111010","111111111111110100","000000000000000010","111111111111101011","111111111111101110","111111111111010111","000000000000000010","000000000000001100","111111111111101111","111111111111101110","000000000000001110","000000000000001000","000000000000000010","111111111111110000","111111111111111100","000000000000000110","000000000000001001","000000000000000100","111111111111011000","000000000000010000","000000000000110011","000000000000000001","111111111111010110"),
("000000000000010101","000000000000001001","000000000000001001","000000000000011111","111111111111010011","000000000000000111","111111111111110110","111111111111011000","111111111111011011","111111111111111100","111111111111111010","000000000000100001","000000000000001100","111111111111001110","000000000000010010","000000000000000010","111111111111110001","111111111111111101","111111111111110001","000000000000001001","000000000000010111","111111111111101101","111111111111011001","111111111111111010","111111111111110101","000000000000110001","111111111111111111","111111111111100101","000000000000000100","000000000000100100","000000000000001010","000000000000101100","111111111111111101","000000000000011010","000000000000100111","111111111111100111","000000000000011000","000000000000001010","111111111111101010","111111111111111101","000000000000001110","000000000000010100","000000000000001100","000000000000001001","111111111111110101","000000000000001011","111111111111111101","000000000000100001","111111111111110111","111111111111101001","111111111111100100","111111111111011100","000000000000000000","000000000000000010","111111111111111101","111111111111111001","111111111111111001","111111111111100011","111111111111010000","000000000000010001","000000000000001001","000000000000011010","111111111111110110","111111111111011111","111111111111111011","111111111111001110","000000000000000000","000000000000011101","000000000000010110","111111111111100100","000000000000100011","000000000000000110","000000000000000001","111111111111101011","000000000000100010","000000000000000100","000000000000010101","111111111111110101","111111111111101001","111111111111101100","111111111111111001","111111111111101101","111111111111100101","111111111111010111","000000000000000111","111111111111011010","000000000000011101","000000000000100011","000000000000011100","000000000000000100","000000000000010101","111111111111100101","111111111111111010","111111111111111110","111111111111010010","000000000000011100","111111111111101001","000000000000010101","000000000000110011","111111111111110011","111111111111111100","111111111111110101","000000000000001100","000000000000010011","111111111111110101","111111111111111011","111111111111111111","000000000000001011","111111111111111101","111111111111100100","111111111111111000","111111111111101100","111111111111111010","111111111111110010","111111111111111111","000000000000000010","111111111111111011","000000000000010100","111111111111100111","111111111111111110","000000000000000000","111111111111101010","000000000000101001","111111111111111010","111111111111111001","000000000000110000","000000000000010001","111111111111001110"),
("000000000000001001","000000000000000001","111111111111101100","000000000000000000","000000000000000001","111111111111111100","000000000000010001","111111111111101001","111111111111011110","000000000000000000","111111111111110001","111111111111111010","111111111111110101","111111111111001110","111111111111111101","000000000000011010","111111111111110011","111111111111111110","000000000000000100","111111111111111101","000000000000010110","111111111111111001","111111111111100101","000000000000000011","000000000000001110","000000000000100110","111111111111111001","111111111111111011","111111111111011101","000000000000101111","000000000000001101","000000000000011010","000000000000000010","000000000000010010","000000000000101011","111111111111111001","000000000000100001","000000000000010001","111111111111111010","000000000000001111","000000000000001111","000000000000101101","111111111111111111","111111111111110011","000000000000000000","111111111111111000","000000000000000000","000000000001000100","111111111111101010","111111111111101101","111111111111010011","111111111111100110","111111111111111100","000000000000001111","000000000000001110","111111111111111000","000000000000010010","111111111111100010","111111111111101001","000000000000001110","000000000000100010","000000000000001000","000000000000000011","111111111111101110","111111111111100100","111111111111101101","000000000000001011","000000000000001100","000000000000011101","000000000000000000","111111111111111101","000000000000001110","000000000000011000","111111111111001110","000000000000110000","000000000000001110","000000000000011000","111111111111100101","000000000000010000","111111111111101101","111111111111010111","000000000000001000","111111111111010100","111111111111010010","000000000000001110","111111111111101110","000000000000010010","000000000000001011","000000000000000001","000000000000001000","111111111111110011","000000000000010000","000000000000010001","111111111111110110","111111111111101000","000000000000101101","111111111111101100","000000000000000111","000000000000000010","111111111111101001","000000000000011100","000000000000001000","000000000000000111","000000000000001111","111111111111111000","000000000000000011","111111111111111111","000000000000000110","111111111111101110","111111111111110101","000000000000000000","000000000000010100","000000000000010011","000000000000000101","111111111111110100","111111111111101011","000000000000010000","000000000000001001","000000000000010001","111111111111111011","000000000000010110","111111111111111111","000000000000000001","000000000000100010","111111111111110001","000000000000011011","000000000000100110","111111111111011000"),
("000000000000000101","000000000000000000","111111111111111001","111111111111101101","000000000000000111","000000000000000011","111111111111101000","111111111111111010","111111111111011010","111111111111101110","111111111111000101","000000000000001011","111111111111110001","111111111111011011","000000000000001011","111111111111101111","111111111111111000","111111111111110110","111111111111010110","111111111111100100","111111111111100111","000000000000001011","000000000000001000","111111111111100001","111111111111111011","111111111111111000","111111111111110010","111111111111001111","111111111111110001","000000000000001000","000000000000000010","000000000000001100","111111111111010111","000000000000110111","000000000000001011","000000000000010101","111111111111111110","000000000000000000","000000000000000010","000000000000000000","000000000000000001","000000000000101001","111111111111101000","000000000000001001","111111111111110100","000000000000001010","111111111111111010","000000000000110110","111111111111110110","000000000000010001","111111111111111000","111111111111111001","000000000000011100","000000000000001111","000000000000000010","111111111111101011","000000000000010101","111111111111101100","111111111111100100","000000000000000000","000000000000011010","111111111111111010","111111111111111111","111111111111111101","000000000000000010","000000000000001001","000000000000001010","000000000000011101","111111111111100011","111111111111101101","000000000000000010","000000000000000100","000000000000101110","111111111111101000","000000000000011101","000000000000100000","111111111111101101","111111111111111001","111111111111110111","111111111111100001","000000000000000001","111111111111011111","111111111111111111","111111111111101000","000000000000000010","111111111111101000","000000000000100111","000000000000101010","000000000000000110","111111111111110001","000000000000010000","111111111111110101","000000000000001010","000000000000000001","111111111110101101","000000000000101000","111111111111111101","000000000000000000","000000000000111000","111111111111010111","000000000000000011","111111111111101101","000000000000001101","000000000000001100","111111111111111010","111111111111011100","111111111111110101","000000000000000000","111111111111111110","000000000000001100","111111111111100000","000000000000000000","000000000000001111","000000000000000111","111111111111101000","111111111111111010","111111111111111110","000000000000010010","000000000000010100","000000000000100001","111111111111111001","000000000000010101","000000000000000011","000000000000010011","000000000000001110","000000000000011101","111111111111111110","111111111111100001"),
("000000000000110000","000000000000000101","111111111111101111","000000000000010001","000000000000001110","111111111111111001","000000000000010101","000000000000000000","111111111111010110","000000000000010000","111111111111010000","000000000000010011","111111111111100010","111111111111011011","111111111111101011","000000000000000011","000000000000001100","111111111111110111","111111111111001001","111111111111101011","111111111111101001","000000000000010001","111111111111111110","111111111111100110","111111111111101010","000000000000011110","111111111111101010","111111111111110001","000000000000010000","000000000000001110","000000000000001111","000000000000000000","111111111111111101","000000000000101001","000000000000001010","000000000000000010","000000000000010010","000000000000001001","111111111111101100","000000000000000011","000000000000011101","000000000000100101","111111111111111001","000000000000100011","111111111111101011","000000000000011000","000000000000000101","000000000001000111","111111111111100111","000000000000011100","111111111111111010","111111111111100010","000000000000011011","000000000000010101","111111111111101110","111111111111001100","000000000000010000","111111111111101110","111111111111011001","111111111111101101","000000000000010100","111111111111110000","111111111111101100","111111111111110110","111111111111110000","111111111111111000","111111111111101001","000000000000010101","111111111111001001","000000000000000001","000000000000011010","111111111111111000","000000000000010101","111111111111101111","000000000000001010","000000000000011000","000000000000001000","111111111111110000","000000000000001001","111111111111101111","000000000000000000","111111111111101110","000000000000001001","111111111111110010","000000000000001011","000000000000001011","000000000000001100","000000000000010101","000000000000001001","111111111111110000","000000000000010111","000000000000001111","000000000000001101","111111111111111001","111111111111011010","000000000000111100","111111111111101100","000000000000000000","000000000000011011","111111111111110001","000000000000010110","000000000000001010","000000000000100100","111111111111110000","111111111111100110","000000000000010011","111111111111100110","000000000000101010","111111111111110001","111111111111101100","111111111111010010","000000000000000000","111111111111111111","111111111111111101","111111111111100111","000000000000010101","000000000000011001","000000000000001001","000000000000000100","000000000000011001","000000000000000011","111111111111110010","111111111111110101","000000000000010000","000000000000010110","000000000000011110","111111111111111000","111111111111011100"),
("000000000000110100","111111111111111101","111111111111101001","111111111111110110","000000000000010100","000000000000000000","000000000000111100","111111111111111111","111111111111100011","000000000000011111","111111111111011001","000000000000011000","111111111111101110","111111111111101001","000000000000001000","000000000000001101","000000000000000110","111111111111111000","111111111111111001","111111111111111001","111111111111011011","000000000000000110","111111111111111110","111111111111010010","111111111111110010","000000000000001110","000000000000000110","111111111111101001","000000000000000111","000000000000000111","000000000000000111","000000000000011001","111111111111110100","000000000000001011","000000000000000000","111111111111100101","111111111111111001","111111111111111101","111111111111011101","111111111111011101","000000000000001001","000000000000011101","111111111111101000","000000000000101000","111111111111010011","000000000000001111","000000000000101000","000000000001001111","111111111111011011","000000000000101011","000000000000000000","111111111111101000","000000000000010001","111111111111111100","111111111111110000","111111111111011001","000000000000010011","111111111111011110","111111111111010010","111111111111110111","000000000000000001","111111111111100101","111111111111110110","000000000000000111","111111111111011000","111111111111110010","111111111111100011","000000000000100001","111111111111001011","111111111111111100","000000000000000011","000000000000010001","000000000000110100","111111111111111111","000000000000011001","000000000000011010","111111111111110000","111111111111110101","000000000000000111","000000000000000010","000000000000000011","111111111111111010","000000000000000111","111111111111111000","000000000000001011","000000000000000001","000000000000001001","000000000000000010","000000000000100001","000000000000000111","111111111111111111","000000000000011000","000000000000011001","000000000000000100","111111111111100110","000000000000000000","111111111111111011","000000000000101111","000000000000101010","111111111111110010","000000000000100111","000000000000011101","000000000000101010","000000000000001001","111111111111110011","000000000000101000","111111111111100001","000000000000100001","111111111111100111","000000000000000011","111111111111011100","000000000000010111","000000000000100011","111111111111001110","111111111111010110","000000000000101000","000000000000001111","000000000000000000","111111111111110100","000000000000001000","000000000000000110","111111111111101100","000000000000000000","000000000000010100","000000000000011101","000000000000010100","000000000000011110","111111111111101100"),
("000000000000100001","000000000000010010","111111111111101100","000000000000000100","000000000000100000","000000000000011011","000000000000010010","000000000000001010","111111111111110001","000000000000010011","000000000000000001","000000000000010111","111111111111110000","111111111111110000","111111111111111111","111111111111110011","111111111111101111","111111111111110010","111111111111110011","111111111111110000","111111111111101110","000000000000010001","000000000000000001","111111111111100000","000000000000000010","000000000000010111","111111111111111100","111111111111101001","000000000000010101","111111111111111100","111111111111101010","000000000000100111","111111111111011000","000000000000110011","111111111111110000","111111111111110101","000000000000000011","111111111111100010","111111111111110111","111111111111101111","000000000000001101","000000000000011010","000000000000010010","000000000000100011","111111111111101000","000000000000000010","000000000000110000","000000000000110001","111111111111111110","000000000000111111","111111111111110111","111111111111010110","000000000000001110","000000000000011001","111111111111111111","111111111111101101","000000000000000101","111111111111110100","111111111111110100","111111111111111000","000000000000011111","111111111111101000","111111111111011001","111111111111111010","111111111111101100","000000000000010100","111111111111100101","000000000000010000","111111111111101101","111111111111111100","000000000000000111","000000000000000100","000000000000100010","000000000000001001","000000000000011111","000000000000001001","111111111111011101","111111111111110010","000000000000010011","111111111111100000","000000000000000100","111111111111010010","000000000000000101","111111111111100101","111111111111101110","000000000000010111","000000000000001010","000000000000010001","000000000000110011","000000000000001100","000000000000100010","000000000000011110","000000000000101100","000000000000100010","111111111111011001","000000000000010010","111111111111110101","000000000000101111","000000000000010111","111111111111110111","000000000000000110","000000000000100101","000000000000100100","111111111111101000","111111111111110110","000000000000000110","111111111111100010","000000000000011111","111111111111110101","111111111111111001","111111111111101100","000000000000000101","000000000000010011","111111111111011100","111111111111100100","000000000000010010","000000000000100101","111111111111111111","000000000000000100","111111111111110111","000000000000001011","000000000000000001","000000000000011011","000000000000100000","000000000000001011","000000000000000111","000000000000011111","111111111111011111"),
("000000000000011111","000000000000001110","111111111111110011","111111111111111100","111111111111110110","000000000000001011","000000000000001110","000000000000001000","111111111111101100","000000000000010111","000000000000010100","000000000000011010","111111111111101011","111111111111110010","111111111111111110","000000000000011001","111111111111101011","111111111111101111","000000000000010000","000000000000000000","111111111111101100","111111111111010001","111111111111011001","111111111111100010","111111111111110101","000000000000001000","111111111111100000","000000000000000110","000000000000001110","111111111111111100","000000000000000000","000000000000001001","111111111111100011","000000000000100110","000000000000000110","111111111111101011","111111111111110010","000000000000000101","000000000000000100","111111111111110100","000000000000000011","000000000000011001","000000000000000000","000000000000011101","111111111111101010","000000000000010000","000000000000000011","000000000000110110","111111111111010100","000000000000010011","111111111111100101","111111111111110110","000000000000101010","000000000000011101","111111111111101101","111111111111001100","000000000000000110","111111111111101010","111111111111101000","111111111111110100","000000000000010101","111111111111101101","111111111111101100","000000000000000010","111111111111111111","000000000000000000","000000000000000101","000000000000010111","111111111111101011","111111111111101110","111111111111110110","000000000000000000","000000000000011101","111111111111110001","000000000000010110","111111111111111011","111111111111101011","111111111111110111","000000000000001011","111111111111011111","111111111111101001","111111111111100111","111111111111101100","111111111111101000","111111111111101000","111111111111100111","000000000000000101","000000000000000110","000000000000001000","000000000000000100","000000000000010111","000000000000001101","000000000000101100","000000000000010011","111111111111011000","000000000000000101","111111111111111100","000000000000011100","000000000000101100","111111111111101100","000000000000010011","000000000000000011","000000000000100001","111111111111100101","000000000000000011","000000000000100010","111111111111101111","000000000000010010","111111111111100101","000000000000000000","111111111111100010","000000000000000100","000000000000011011","111111111111111110","111111111111000110","000000000000010110","000000000000000101","000000000000001110","111111111111110000","000000000000011010","000000000000001110","111111111111110101","000000000000001111","000000000000011100","000000000000011001","111111111111111110","000000000000010101","111111111111100000"),
("000000000000010010","111111111111111101","111111111111101001","111111111111110111","111111111111101011","111111111111111111","000000000000100000","111111111111111001","000000000000001001","111111111111111001","111111111111111100","111111111111110111","000000000000001001","111111111111101110","000000000000010001","000000000000011100","000000000000010100","000000000000001000","000000000000011111","000000000000001100","111111111111111001","111111111111101110","111111111111111011","111111111111100010","111111111111101100","000000000000001010","111111111111100110","000000000000001111","000000000000000100","000000000000010010","000000000000000100","111111111111111100","111111111111111010","000000000000000100","000000000000011001","111111111111101000","000000000000001101","000000000000001111","111111111111111010","111111111111110101","111111111111110001","000000000000001011","000000000000001110","000000000000000010","111111111111100111","111111111111110111","000000000000000011","111111111111101101","111111111111011110","000000000000000010","111111111111110110","111111111111111110","111111111111111000","000000000000011110","111111111111110110","111111111111011010","111111111111011101","111111111111101011","111111111111010110","111111111111111000","111111111111110010","111111111111111101","000000000000000111","000000000000000011","000000000000010100","111111111111101010","111111111111111011","111111111111111111","000000000000000000","000000000000000111","111111111111111111","000000000000011000","111111111111110110","000000000000000011","111111111111110100","111111111111111111","000000000000000000","000000000000001101","111111111111111000","000000000000001001","111111111111111000","111111111111101000","000000000000010010","111111111111101011","000000000000001001","111111111111111011","111111111111111001","111111111111111111","111111111111111100","111111111111111111","111111111111101110","000000000000001101","111111111111101110","000000000000001110","111111111111101000","000000000000001101","000000000000010010","000000000000000011","111111111111110000","111111111111101101","000000000000100010","111111111111110100","000000000000001100","000000000000000100","111111111111111010","000000000000010100","111111111111101010","000000000000000000","000000000000001010","000000000000001001","111111111111011110","000000000000001110","000000000000010001","111111111111101110","000000000000011001","000000000000100111","000000000000010001","111111111111110111","000000000000000001","000000000000000111","000000000000000000","111111111111110111","000000000000001011","000000000000100001","111111111111111011","000000000000000000","000000000000100100","111111111111110101"),
("111111111111101100","111111111111101011","111111111111101101","000000000000010111","000000000000001010","111111111111111000","000000000000100000","000000000000010011","000000000000011110","111111111111110110","000000000000100001","111111111111110100","000000000000011011","111111111111111001","000000000000001110","000000000000011111","000000000000100010","000000000000001101","000000000000001001","000000000000010011","000000000000000110","111111111111111011","111111111111111000","000000000000001000","111111111111101000","000000000000011001","111111111111111011","000000000000001100","000000000000010101","111111111111111110","000000000000000000","000000000000001110","000000000000011001","000000000000001000","000000000000000011","000000000000001011","000000000000001001","000000000000000001","000000000000000011","111111111111101100","111111111111111100","111111111111101101","000000000000011100","000000000000011100","111111111111111111","000000000000010101","111111111111101010","000000000000001001","000000000000000100","000000000000010110","000000000000011010","111111111111111110","111111111111110101","000000000000001110","111111111111101110","111111111111101001","111111111111101001","000000000000010001","111111111111110100","111111111111110001","111111111111111011","000000000000001101","000000000000000000","111111111111101111","111111111111110110","111111111111100100","111111111111111011","111111111111110000","000000000000011000","000000000000001000","000000000000010010","000000000000001010","000000000000000101","111111111111101110","111111111111111110","111111111111111110","000000000000010010","111111111111110010","111111111111111100","111111111111110111","000000000000000100","000000000000010101","111111111111111101","111111111111101011","000000000000010010","111111111111111000","000000000000000111","111111111111101011","000000000000000001","111111111111101001","000000000000001001","111111111111101100","111111111111110011","111111111111111011","000000000000000000","000000000000000010","000000000000000101","111111111111111000","111111111111101111","000000000000000111","000000000000001100","111111111111110110","000000000000010001","000000000000000100","000000000000000110","000000000000010010","000000000000000101","000000000000010011","111111111111101111","000000000000001111","111111111111011101","000000000000000111","000000000000000111","111111111111101110","000000000000010111","000000000000010010","111111111111110111","000000000000010001","000000000000000100","000000000000001001","111111111111110100","000000000000000010","000000000000001010","111111111111110010","111111111111111001","000000000000000000","000000000000010110","111111111111110101"),
("111111111111111101","000000000000001101","000000000000000001","000000000000010010","111111111111111010","000000000000000000","000000000000000010","111111111111110101","000000000000000110","000000000000001110","111111111111110100","000000000000001100","000000000000000110","000000000000000100","000000000000001100","000000000000000111","000000000000000100","111111111111110111","000000000000001010","111111111111110011","111111111111111000","111111111111101110","000000000000000000","111111111111101100","000000000000001000","000000000000000101","000000000000000000","111111111111110101","000000000000001101","111111111111110001","111111111111111000","111111111111101110","000000000000000100","000000000000000011","000000000000000100","000000000000000010","000000000000000110","000000000000010100","111111111111110011","000000000000010000","111111111111110010","111111111111110110","111111111111111011","111111111111110100","111111111111110000","000000000000000100","000000000000010010","000000000000010011","111111111111111011","000000000000000010","000000000000000111","111111111111111001","111111111111101111","000000000000000100","111111111111111110","111111111111110011","000000000000000000","111111111111110101","000000000000000000","111111111111111010","111111111111110000","111111111111110001","000000000000000100","000000000000000000","000000000000010010","111111111111111011","111111111111101111","000000000000001000","000000000000001100","000000000000010011","111111111111111101","111111111111110000","000000000000001000","000000000000010000","111111111111111001","000000000000000001","111111111111111100","111111111111101101","000000000000001110","111111111111111001","111111111111111100","111111111111110010","111111111111101110","000000000000001000","111111111111111111","111111111111110010","000000000000001111","000000000000001010","000000000000000101","111111111111111110","000000000000000011","111111111111111100","111111111111111011","111111111111110000","111111111111110101","111111111111101110","111111111111110101","000000000000001000","000000000000001011","111111111111111111","111111111111111000","111111111111111111","000000000000000001","111111111111101110","111111111111110111","111111111111101101","000000000000000101","000000000000010010","000000000000001011","000000000000001110","111111111111110100","111111111111110110","111111111111111110","000000000000000101","111111111111110111","000000000000000101","000000000000000000","000000000000000110","111111111111111001","111111111111111000","000000000000000010","111111111111110100","000000000000000011","000000000000010001","111111111111111001","000000000000001001","111111111111101110","111111111111101100"),
("000000000000001010","111111111111110000","000000000000001000","000000000000010011","000000000000001001","000000000000001110","111111111111110100","000000000000000011","000000000000000101","000000000000001001","111111111111110001","111111111111101100","000000000000010010","000000000000001110","111111111111111010","111111111111101110","000000000000001001","111111111111110010","111111111111110111","000000000000010010","000000000000010001","000000000000000011","000000000000001001","000000000000000100","111111111111110101","000000000000010001","000000000000000100","111111111111111010","111111111111111110","000000000000001101","111111111111101110","000000000000000000","000000000000000010","000000000000010001","111111111111111110","000000000000000011","000000000000010010","111111111111101100","111111111111101101","111111111111110101","111111111111110111","111111111111111001","111111111111110011","000000000000001111","000000000000000100","000000000000001010","111111111111110110","111111111111111111","111111111111111100","000000000000010011","111111111111110101","111111111111111011","000000000000010001","111111111111111001","000000000000000011","111111111111111101","000000000000000111","111111111111101100","000000000000001000","000000000000000101","111111111111110000","111111111111111101","111111111111111110","000000000000000100","000000000000010100","111111111111110011","111111111111111101","111111111111110001","000000000000000110","000000000000000010","111111111111101110","000000000000000110","111111111111110100","111111111111110101","000000000000000001","000000000000010100","000000000000001001","000000000000000010","111111111111111101","111111111111111001","000000000000001001","000000000000000100","000000000000000101","111111111111111110","111111111111111101","000000000000010100","000000000000000010","111111111111101100","000000000000000100","000000000000000110","000000000000001010","111111111111111111","000000000000000000","111111111111110010","111111111111111010","111111111111111001","000000000000001111","000000000000001011","111111111111111010","111111111111101101","111111111111111100","111111111111111011","111111111111111001","000000000000001111","000000000000000000","000000000000000011","111111111111110101","111111111111111011","000000000000010011","000000000000010011","111111111111101100","000000000000001011","000000000000000110","111111111111101101","111111111111111011","111111111111111101","111111111111110000","111111111111111100","111111111111101110","111111111111111111","111111111111110110","111111111111111100","000000000000000110","111111111111101101","000000000000010100","000000000000001111","111111111111111011","000000000000010001"),
("000000000000010000","000000000000010000","111111111111111001","111111111111110100","111111111111110011","000000000000000101","111111111111110010","000000000000001111","000000000000000010","000000000000001101","000000000000000001","000000000000001110","000000000000010010","000000000000001101","000000000000000000","000000000000000011","111111111111110100","000000000000000010","111111111111111110","000000000000000000","111111111111111100","111111111111101111","000000000000001011","000000000000010001","111111111111110001","111111111111110111","111111111111101110","000000000000001000","111111111111110100","000000000000010011","000000000000000000","000000000000000000","000000000000001111","111111111111111001","111111111111111001","111111111111111011","111111111111111101","111111111111111111","111111111111111010","111111111111111000","000000000000001011","000000000000010100","000000000000001111","000000000000000100","000000000000001110","111111111111110111","111111111111111101","000000000000000001","000000000000000110","111111111111111111","111111111111110001","000000000000010001","000000000000000010","111111111111111011","000000000000000000","111111111111111010","111111111111111011","000000000000001100","111111111111111111","111111111111111011","111111111111111110","000000000000000110","111111111111101101","000000000000001111","111111111111101101","111111111111111001","000000000000010001","000000000000001101","111111111111110010","000000000000010011","111111111111101110","000000000000000100","000000000000000111","111111111111110111","000000000000000111","000000000000001011","111111111111110011","111111111111110110","000000000000001011","111111111111110001","000000000000000111","000000000000010001","111111111111110001","000000000000000000","111111111111111101","111111111111101111","111111111111111001","111111111111110001","000000000000000000","000000000000000000","111111111111110110","111111111111111110","000000000000000111","000000000000010000","111111111111111000","000000000000001111","111111111111110000","111111111111110100","111111111111111011","111111111111111001","000000000000001001","111111111111111101","111111111111110100","111111111111111011","111111111111111100","111111111111101111","000000000000001011","000000000000001000","111111111111111100","000000000000010100","000000000000001110","111111111111110100","111111111111111101","000000000000010100","111111111111111001","000000000000010011","111111111111111100","000000000000001000","111111111111111011","111111111111111001","111111111111101110","000000000000010010","111111111111111001","111111111111110101","000000000000010010","111111111111101100","000000000000000011","000000000000010001"),
("000000000000001101","111111111111101110","111111111111110010","111111111111110010","000000000000010000","000000000000000101","000000000000001111","000000000000000110","000000000000001011","111111111111111010","111111111111111011","111111111111101110","111111111111111011","111111111111111100","111111111111110010","111111111111111111","111111111111111001","000000000000001010","111111111111101111","111111111111111000","111111111111110101","000000000000000000","000000000000001011","000000000000001000","000000000000001010","111111111111111000","000000000000000101","000000000000001000","111111111111110101","111111111111110101","000000000000000000","111111111111110111","000000000000000100","111111111111110110","000000000000000100","111111111111111110","000000000000001000","000000000000000001","111111111111110100","000000000000001100","111111111111110111","000000000000000110","000000000000010011","111111111111111010","111111111111110011","000000000000010010","000000000000010100","111111111111111000","000000000000010001","111111111111110111","000000000000000000","000000000000000101","111111111111110000","000000000000010010","111111111111111000","000000000000001010","111111111111110001","000000000000000010","111111111111101101","111111111111111001","000000000000000000","000000000000000111","000000000000000111","000000000000000001","111111111111111100","000000000000001111","111111111111101110","111111111111101110","111111111111110010","000000000000000101","000000000000000111","111111111111110001","000000000000001110","111111111111111101","000000000000000000","000000000000001001","000000000000010000","000000000000001001","000000000000000000","111111111111110111","111111111111110010","000000000000000110","000000000000010011","000000000000000111","111111111111101101","111111111111111011","000000000000000111","000000000000000111","111111111111111110","111111111111110100","000000000000000000","000000000000000011","111111111111111001","111111111111110100","000000000000010000","000000000000001000","111111111111101110","111111111111110010","111111111111101101","000000000000001100","000000000000001011","000000000000000001","000000000000000110","000000000000000001","111111111111110111","111111111111101101","000000000000000001","111111111111111110","111111111111111011","111111111111110111","111111111111111000","111111111111110010","111111111111101111","000000000000010011","111111111111111000","111111111111111110","000000000000000010","111111111111111011","000000000000001100","111111111111110110","111111111111110010","111111111111101101","000000000000010011","000000000000000111","111111111111110111","000000000000001101","000000000000010001","000000000000010001"),
("111111111111100111","000000000000010011","111111111111101010","000000000000011100","000000000000011110","111111111111110000","111111111111101010","000000000000000110","000000000000010010","000000000000000001","000000000000100110","111111111111111111","000000000000011000","000000000000010000","000000000000010010","111111111111110000","111111111111100010","000000000000011100","000000000000010001","111111111111111011","000000000000010011","000000000000000000","000000000000000001","000000000000011100","000000000000000101","000000000000010000","000000000000010010","000000000000001100","000000000000001101","000000000000010010","000000000000101000","111111111111011111","111111111111111000","000000000000001101","000000000000101000","000000000000000110","111111111111111001","000000000000100100","111111111111111111","000000000000001100","000000000000010010","000000000000010001","111111111111111011","000000000000011101","111111111111011100","000000000000101110","111111111111010111","000000000000001011","111111111111010101","111111111111111001","000000000000000000","111111111111010111","111111111111111111","000000000000000101","000000000000011111","000000000000001100","111111111111101110","111111111111110001","111111111111110011","000000000000000111","111111111111011001","000000000000101000","000000000000000101","000000000000000101","000000000000001100","111111111111100100","111111111111110011","111111111111100110","000000000000000111","000000000000000100","000000000000100000","000000000000011101","111111111111010100","000000000000011101","000000000000010000","111111111111100000","111111111111101010","000000000000001000","000000000000000110","111111111111011110","000000000000010010","111111111111101110","000000000000010010","000000000000010011","000000000000011010","111111111111111100","111111111111110000","111111111111110101","111111111111101101","000000000000100101","000000000000100001","111111111111101101","111111111111110111","000000000000011111","111111111111111111","111111111111100110","000000000000001101","000000000000000000","111111111111110010","111111111111101110","111111111111100101","000000000000001100","111111111111101110","000000000000010100","000000000000011110","111111111111110010","000000000000000110","111111111111111010","000000000000001101","000000000000000101","000000000000100010","000000000000001010","111111111111111011","111111111111011101","000000000000001101","111111111111110110","111111111111100001","000000000000010010","000000000000011110","000000000000101010","000000000000000100","111111111111111001","000000000000001001","000000000000000001","111111111111011010","111111111111101011","111111111111110111","000000000000101000"),
("000000000000001101","111111111111111101","111111111111110000","000000000000000011","111111111111101100","111111111111110100","000000000000011000","000000000000000011","000000000000000100","000000000000000110","111111111111111001","111111111111101110","000000000000000111","000000000000001110","111111111111101010","111111111111110110","111111111111100000","000000000000010010","000000000000011000","000000000000001001","000000000000010110","111111111111111100","111111111111111010","111111111111111011","111111111111111000","000000000000000000","000000000000000101","000000000000000010","111111111111111100","111111111111111000","111111111111101001","000000000000011101","111111111111111101","000000000000100110","000000000000001010","000000000000011101","000000000000000101","111111111111110001","111111111111011010","111111111111100011","111111111111111100","000000000000100100","000000000000100101","000000000000000000","111111111111101111","111111111111110001","000000000000100110","000000000000010000","111111111111111000","111111111111100110","000000000000010001","111111111111100010","000000000000100011","111111111111110110","000000000000001010","111111111111110110","111111111111011111","111111111111111011","000000000000010000","000000000000000000","000000000000010111","000000000000001000","111111111111111101","111111111111101010","000000000000010100","111111111111110110","000000000000011100","000000000000100000","000000000000001111","000000000000010000","000000000000001111","000000000000001010","000000000000101000","111111111111110000","000000000000001011","000000000000000100","111111111111011001","000000000000010000","111111111111101100","111111111111010101","111111111111100100","111111111111100101","111111111111110010","000000000000001001","111111111111110011","000000000000000001","000000000000000011","000000000000000110","000000000000011010","000000000000000010","111111111111110110","000000000000011001","000000000000110011","000000000000010111","111111111111111111","000000000000001101","111111111111101010","000000000000001111","111111111111111110","111111111111101000","000000000000011000","111111111111101011","000000000000011010","000000000000011100","111111111111111001","000000000000001010","111111111111101001","000000000000000100","111111111111101100","111111111111110110","111111111111100111","111111111111110100","111111111111110010","111111111111111110","111111111111010000","000000000000100000","000000000000000111","000000000000001010","111111111111101000","000000000000010000","000000000000000110","111111111111110111","000000000000011110","000000000000000001","000000000000000100","000000000000010101","111111111111110001","111111111111110000"),
("000000000000100101","111111111111111010","000000000000010000","111111111111100110","111111111111110001","111111111111100111","111111111111111011","111111111111111000","111111111111110011","111111111111111000","000000000000000110","111111111111111001","000000000000010101","000000000000001010","111111111111101101","111111111111011100","111111111111100110","000000000000001010","000000000000000101","111111111111110011","111111111111111100","000000000000001000","111111111111010011","000000000000001001","000000000000011000","111111111111111110","111111111111101111","111111111111101111","111111111111101011","000000000000000011","000000000000000110","111111111111111111","111111111111111011","000000000000011000","000000000000010110","111111111111110001","000000000000100011","111111111111111101","111111111111111110","000000000000011001","111111111111110010","000000000000001000","000000000000000000","000000000000000101","000000000000000100","000000000000000000","000000000000001011","000000000000010000","000000000000001101","111111111111100100","111111111111010111","111111111111110000","000000000000011000","111111111111110010","111111111111111101","111111111111101110","111111111111110110","111111111111110011","111111111111101101","111111111111111100","000000000000100010","000000000000000010","111111111111110100","111111111111011011","111111111111111100","000000000000100011","000000000000101101","111111111111111010","111111111111100011","000000000000010111","111111111111100011","111111111111101011","000000000000100110","000000000000000110","000000000000101001","000000000000000110","000000000000100011","000000000000010101","111111111111111010","111111111111101010","000000000000001110","000000000000001010","111111111111011110","111111111111111101","000000000000001000","111111111111101110","000000000000000000","000000000000110010","000000000000000000","000000000000011011","000000000000010000","111111111111101010","000000000000100110","111111111111111101","111111111111100011","000000000000010010","000000000000000011","000000000000001111","000000000000101010","111111111111010111","000000000000100001","111111111111110100","000000000000000000","000000000000000110","000000000000000011","111111111111110010","000000000000000100","000000000000011111","000000000000010000","111111111111111010","111111111111111110","111111111111101011","111111111111110111","111111111111111001","111111111111101010","111111111111011111","000000000000000101","111111111111111100","111111111111110100","000000000000001100","000000000000110011","000000000000000010","000000000000010010","000000000000000000","111111111111100010","000000000000010010","000000000000001001","000000000000001010"),
("111111111111101001","000000000000010111","111111111111110000","111111111111101001","000000000000010111","111111111111111010","111111111111110011","000000000000011011","000000000000001101","000000000000000011","111111111111110001","111111111111111000","111111111111111110","111111111111100110","000000000000011100","111111111111101101","000000000000011010","111111111111011001","000000000000000111","000000000000001011","111111111111100011","111111111111111010","111111111111100001","111111111111110011","000000000000000000","000000000000011111","111111111111011100","111111111111110011","000000000000010100","000000000000010101","111111111111011111","000000000000000001","000000000000001110","111111111111101110","000000000000000001","111111111111110101","000000000000001100","111111111111101010","000000000000001011","000000000000001100","111111111111111001","111111111111110011","000000000000000000","000000000000001001","000000000000011101","111111111111111011","000000000000101010","000000000000000001","111111111111111110","000000000000010010","000000000000001001","111111111111100001","111111111111111101","111111111111111100","000000000000001010","111111111111011001","000000000000000110","000000000000010010","111111111111011011","000000000000000010","000000000000011110","000000000000001001","111111111111101010","111111111111110010","111111111111100000","111111111111100101","000000000000000010","000000000000100001","111111111111100100","111111111111110011","000000000000001011","000000000000010111","000000000000000000","111111111111101011","000000000000011110","000000000000001100","000000000000000110","000000000000001110","000000000000010111","111111111111111010","000000000000001100","000000000000010100","111111111111111100","111111111111110001","111111111111111100","111111111111111000","111111111111011011","000000000000011101","000000000000100100","000000000000010010","111111111111100100","000000000000000011","000000000000001101","111111111111111011","111111111111011000","000000000000001011","000000000000001101","000000000000001111","000000000000001110","111111111111101011","000000000000010000","000000000000000010","000000000000011111","111111111111101110","111111111111101111","000000000000001011","111111111111100110","000000000000010011","111111111111100110","000000000000000010","111111111111010101","000000000000000000","000000000000010010","000000000000000011","111111111111110010","111111111111111101","000000000000001100","111111111111101111","111111111111101011","000000000000010001","111111111111111101","111111111111110000","111111111111111110","000000000000000110","000000000000000110","111111111111110011","111111111111110101","111111111111011101"),
("111111111111100010","000000000000000100","111111111111110011","000000000000010000","111111111111110111","000000000000011001","111111111111111111","111111111111111001","000000000000000000","000000000000000000","000000000000000100","000000000000000001","000000000000000000","111111111111111000","000000000000110000","000000000000001000","000000000000001000","111111111111111001","000000000000001011","111111111111110110","111111111111100011","111111111111111010","111111111111010011","111111111111101101","111111111111110000","000000000000011010","111111111111100011","111111111111110011","000000000000101100","000000000000000111","000000000000000010","000000000000100100","111111111111111010","111111111111101111","111111111111101011","111111111111111110","111111111111100111","111111111111100111","000000000000000110","000000000000001110","000000000000000011","111111111111100100","000000000000100001","000000000000000001","111111111111101110","111111111111101000","000000000000110000","000000000000000100","000000000000000110","000000000000100001","111111111111100001","111111111111111001","111111111111100001","111111111111100011","000000000000001011","111111111111100011","111111111111101110","000000000000000101","111111111111001111","111111111111110100","111111111111110111","000000000000000100","000000000000001000","000000000000000010","111111111111110011","111111111111011010","000000000000000111","000000000000100110","111111111111101111","111111111111111101","000000000000101100","000000000000000111","111111111111110000","111111111111110101","000000000000101000","000000000000001111","111111111111100100","000000000000010110","000000000000000011","111111111111100011","111111111111110001","000000000000000001","000000000000000010","111111111111100001","111111111111111110","111111111111011001","111111111111100011","000000000000001110","000000000000100010","111111111111110100","111111111111101010","000000000000001110","000000000000011011","000000000000010001","111111111111101100","111111111111101110","000000000000001101","000000000000011111","111111111111111110","111111111111100110","111111111111111110","000000000000011001","000000000000001100","111111111111101101","111111111111110001","000000000000001011","111111111111100001","000000000000010010","111111111111101011","111111111111101111","111111111111011000","111111111111111110","000000000000101010","111111111111110100","111111111111011110","000000000000010010","000000000000110000","111111111111111111","000000000000000010","111111111111111100","111111111111111100","000000000000000100","000000000000000111","111111111111111000","000000000000000110","111111111111111110","111111111111101110","111111111111101000"),
("000000000000000000","000000000000011101","111111111111001100","111111111111111011","111111111111101011","111111111111111110","111111111111101100","111111111111111100","000000000000000100","000000000000100101","111111111111110111","111111111111111111","000000000000001000","000000000000011000","000000000000100001","111111111111111011","000000000000000110","111111111111011001","111111111111111000","000000000000001100","111111111111101101","111111111111101100","111111111111101100","111111111111111001","000000000000000001","000000000000000111","111111111111011011","000000000000010011","000000000000001011","000000000000010100","111111111111110000","000000000000100110","000000000000001000","000000000000000000","111111111111100001","111111111111110011","111111111111101111","000000000000001000","000000000000000000","000000000000000011","111111111111101101","111111111111101011","000000000000010101","000000000000001010","000000000000000010","111111111111101110","000000000000101010","111111111111111111","111111111111110100","000000000000011110","111111111111110100","111111111111110111","111111111111110110","000000000000010010","000000000000001000","111111111111011111","111111111111110101","111111111111101010","111111111111110001","111111111111110000","000000000000011011","000000000000001001","111111111111110011","000000000000001000","000000000000000000","111111111111110001","000000000000001100","000000000000001110","000000000000000100","111111111111100100","000000000000110000","111111111111110111","000000000000000110","111111111111110101","000000000000100111","000000000000001010","111111111111100110","000000000000100111","111111111111111111","111111111111101101","111111111111111010","111111111111110110","000000000000011000","111111111111110011","000000000000000011","111111111111010110","111111111111011010","000000000000101110","000000000000101101","000000000000000010","000000000000001010","000000000000000000","000000000000000111","000000000000010010","111111111111000010","111111111111110000","000000000000011010","000000000000101011","111111111111101001","111111111111111000","000000000000001001","111111111111110000","000000000000011100","000000000000001011","111111111111111000","111111111111110011","111111111111010010","000000000000000100","111111111111010110","111111111111111110","111111111111100110","111111111111101101","000000000000001110","000000000000000010","111111111111111011","000000000000001100","000000000000100101","000000000000000000","111111111111111000","000000000000100101","000000000000010011","111111111111101010","111111111111110110","111111111111111111","000000000000010011","111111111111110111","000000000000001000","111111111111010011"),
("111111111111110111","000000000000110000","111111111111000111","000000000000010000","111111111111110010","000000000000001010","000000000000000100","000000000000011111","111111111111100001","000000000000000110","000000000000001010","111111111111111111","000000000000001000","000000000000000011","000000000000000001","000000000000001110","000000000000000001","111111111111100110","111111111111111000","000000000000011001","111111111111011100","111111111111101101","111111111111100101","111111111111101011","111111111111101001","000000000000010100","111111111111011001","000000000000100111","000000000000000000","111111111111101110","000000000000000111","000000000000011101","000000000000101010","111111111111101100","111111111111110001","111111111111101000","111111111111111111","111111111111111010","111111111111011110","111111111111110000","111111111111111000","111111111111011101","000000000000010010","111111111111111101","000000000000010001","111111111111001110","000000000000110011","111111111111110111","000000000000000111","000000000000001011","000000000000000011","111111111111110011","111111111111110100","000000000000010000","000000000000011010","111111111111011111","111111111111110001","000000000000000010","111111111111110111","000000000000000000","000000000000001011","000000000000001011","000000000000011011","111111111111101000","111111111111011011","111111111111011110","111111111111001100","000000000000100010","000000000000010101","111111111111110100","000000000000100101","000000000000001101","000000000000000101","111111111111111011","000000000000100000","000000000000100011","111111111111101111","000000000000011111","111111111111100010","111111111111110110","111111111111101010","000000000000001001","000000000000001110","111111111111010100","000000000000011010","111111111111010010","111111111111100100","000000000000001101","000000000000001101","000000000000011100","111111111111101000","000000000000011001","000000000000010011","111111111111110110","111111111110110011","111111111111110100","000000000000100100","000000000000110100","111111111111010000","111111111111111111","000000000000000100","000000000000001111","000000000000010011","000000000000000101","111111111111010110","111111111111111011","111111111111001111","000000000000011110","111111111111100100","111111111111111011","111111111110110001","111111111111101100","000000000000100000","000000000000011011","111111111111000111","000000000000110001","000000000001000010","000000000000001100","111111111111111010","000000000000100100","111111111111110111","111111111111011111","111111111111100001","111111111111100011","111111111111101100","000000000000001101","111111111111101100","111111111111100110"),
("000000000000000011","000000000000011101","111111111111000111","000000000000100100","111111111111100111","111111111111111101","000000000000011001","000000000000001101","000000000000000000","111111111111111001","000000000000010101","111111111111111011","000000000000000011","000000000000000111","000000000000001000","000000000000000011","000000000000000111","000000000000011001","000000000000011001","000000000000100000","111111111111010111","111111111111111100","111111111111101000","111111111111111100","111111111111100010","000000000000101011","111111111111010001","000000000000011000","111111111111111111","111111111111101111","000000000000001110","000000000000010100","000000000000110000","111111111111110000","000000000000001000","111111111111001100","000000000000100010","000000000000010001","111111111111011110","111111111111100100","000000000000010010","111111111111100100","000000000000001100","000000000000010110","111111111111111001","111111111111100011","000000000000010101","000000000000010001","111111111111011010","000000000000011111","111111111111100111","111111111111101000","000000000000000000","000000000000110111","000000000000010110","111111111111100010","111111111111111010","111111111111101101","111111111111110001","000000000000001111","000000000000010110","000000000000011011","000000000000100000","111111111111011101","111111111111101001","111111111111011101","111111111111100010","000000000000010010","000000000000000000","111111111111101101","000000000000110110","000000000000010101","111111111111111001","111111111111101100","111111111111111110","000000000000100110","000000000000000000","000000000000100010","111111111111010011","111111111111100110","111111111111110001","000000000000001010","111111111111111000","111111111111101000","111111111111110000","111111111111001111","111111111111011000","000000000000000011","111111111111110001","000000000000000110","111111111111100111","000000000000000010","000000000000100011","000000000000000100","111111111110111111","000000000000000110","000000000000001011","000000000000101111","111111111111011000","111111111111101000","000000000000001010","000000000000000011","000000000000010001","000000000000000101","111111111111111000","000000000000011001","111111111110111010","000000000000100110","111111111111011010","111111111111111010","111111111111010101","111111111111100100","000000000000011010","111111111111101010","111111111111000001","000000000000110011","000000000000100101","000000000000010110","111111111111010110","000000000000111101","000000000000101010","000000000000001001","000000000000010001","111111111111111000","000000000000011110","111111111111110110","000000000000011010","111111111111100001"),
("111111111111100110","000000000000000011","111111111111001101","000000000000011000","111111111111111010","000000000000010010","000000000000000011","000000000000101010","000000000000000111","000000000000000111","000000000000001100","000000000000011101","000000000000000000","111111111111101110","111111111111111111","000000000000011000","000000000000001010","000000000000010001","111111111111111010","000000000000001111","111111111110110100","000000000000000111","111111111111011101","111111111111100010","111111111111101111","000000000000011011","111111111111000110","000000000000010010","000000000000001100","111111111111011000","111111111111101101","000000000000000000","000000000000101011","111111111111101101","111111111111111010","111111111111100000","111111111111111100","000000000000011010","111111111111010011","111111111111110111","000000000000001110","111111111111100011","111111111111111110","111111111111101100","111111111111111001","111111111111110100","000000000000011011","000000000000001000","000000000000001011","000000000000010101","111111111111111010","111111111111101100","000000000000000010","000000000000011001","000000000000010100","111111111111011110","111111111111110111","000000000000011001","111111111111100111","111111111111101100","111111111111111111","000000000000010100","000000000000011001","111111111111010010","111111111111011001","111111111111011110","111111111111100010","000000000000001000","111111111111011110","111111111111111000","000000000000001011","000000000000011100","000000000000000101","111111111111111011","000000000000001010","000000000000101110","111111111111111101","000000000000011110","111111111111101010","000000000000000011","111111111111001001","000000000000100011","000000000000010000","111111111111110010","000000000000001100","111111111111100110","111111111111111001","000000000000000011","111111111111101111","000000000000001110","111111111111011001","111111111111111010","000000000000001100","111111111111111000","111111111111001110","111111111111111100","000000000000011100","000000000000100110","111111111111011001","000000000000001100","111111111111111111","000000000000001110","111111111111111000","000000000000000001","111111111111101001","000000000000001101","111111111111010111","000000000000001111","111111111111010000","111111111111011111","111111111111001001","111111111111100101","111111111111111101","111111111111111010","111111111110100101","000000000000010001","000000000000101111","000000000000001101","111111111111011110","000000000000011101","000000000000011110","111111111111100111","000000000000001010","111111111111110111","111111111111111100","111111111111101000","111111111111111100","111111111111010100"),
("000000000000000000","000000000000001111","111111111111001101","000000000000011001","111111111111101010","000000000000001100","000000000000011001","000000000000011111","000000000000010100","000000000000001100","111111111111110011","111111111111111001","111111111111110100","111111111111100011","000000000000000111","000000000000001011","000000000000000000","000000000000001010","111111111111110100","000000000000101010","111111111110110011","111111111111101101","000000000000000000","111111111111100001","111111111111100111","000000000000010100","111111111111010000","000000000000001100","000000000000011100","111111111111110111","111111111111101110","000000000000000000","000000000000110100","111111111111011011","000000000000000101","111111111111101001","000000000000000111","000000000000001001","111111111111111110","111111111111110101","111111111111111011","111111111111010010","111111111111110101","111111111111110010","000000000000101011","111111111111100100","000000000000101000","111111111111111001","111111111111110011","000000000000010001","111111111111111011","000000000000010000","111111111111100011","000000000000000010","000000000000100100","111111111111100110","111111111111101101","000000000000000110","111111111111101111","000000000000010010","000000000000100000","000000000000011001","000000000000000001","111111111111110000","111111111111010010","111111111111010110","111111111111101000","000000000000001111","111111111111011010","111111111111011101","000000000000010100","000000000000001010","111111111111111000","000000000000010001","111111111111111011","000000000000011110","000000000000000010","000000000000101010","111111111111110011","111111111111110101","111111111111100111","000000000000101011","000000000000010000","111111111111111101","000000000000001101","111111111111100110","111111111111010110","000000000000011011","000000000000001101","000000000000010100","111111111111100000","000000000000001100","000000000000110101","111111111111100111","111111111111000100","000000000000000000","000000000000010110","000000000000011111","111111111111111111","111111111111110001","000000000000010101","000000000000101000","111111111111111110","000000000000000000","111111111111001101","000000000000010010","111111111110110101","000000000000001000","111111111111011100","000000000000001000","111111111111010100","111111111111110110","000000000000001011","111111111111101111","111111111110110010","000000000000011011","000000000000011100","000000000000010101","111111111111100010","000000000000011111","000000000000010011","111111111111111010","000000000000001110","111111111111000101","000000000000001101","111111111111011100","000000000000100001","111111111111100000"),
("111111111111110001","000000000000111010","111111111111001001","000000000000100000","111111111110111111","000000000000010111","000000000000000011","000000000000100000","111111111111110111","000000000000001110","111111111111111111","000000000000001010","111111111111101110","111111111111110111","000000000000011101","000000000000001100","000000000000000100","000000000000010111","111111111111111001","000000000000000110","111111111111101001","111111111111011110","111111111111111000","111111111111101110","111111111111111111","000000000000001101","111111111111010011","000000000000010000","000000000000010010","111111111111111011","111111111111110100","000000000000101001","000000000000001011","111111111111100110","000000000000010011","111111111111010011","000000000000010000","000000000000001001","000000000000010011","000000000000001100","000000000000011011","111111111111100001","000000000000000001","000000000000000010","000000000000010100","111111111111111000","000000000000011110","000000000000000010","111111111111101110","111111111111111101","000000000000001010","000000000000001000","111111111111111000","000000000000000000","000000000000001010","111111111111010100","111111111111111001","000000000000001000","111111111111101000","111111111111111011","000000000000000110","000000000000110011","000000000000011010","111111111111011011","111111111111101110","111111111111110001","111111111111110010","000000000000100101","111111111111110011","111111111111100101","000000000000100100","000000000000101101","000000000000001000","000000000000000100","000000000000010100","000000000000011001","000000000000001010","000000000000100011","111111111111101000","111111111111011101","111111111111010001","111111111111111100","000000000000001101","111111111111100101","000000000000010110","111111111111110000","111111111111100011","000000000000001111","111111111111101010","111111111111111000","000000000000011000","111111111111111001","000000000000010110","111111111111111000","111111111110111110","000000000000000001","000000000000011110","000000000000010111","111111111111110100","111111111111111010","111111111111111100","000000000000101101","111111111111110110","000000000000010110","111111111111101010","000000000000010011","111111111110101001","000000000000100001","111111111111010110","111111111111101100","111111111111011001","111111111111110001","000000000000011110","000000000000010100","111111111110100000","000000000000001111","000000000000101011","000000000000010110","111111111111011111","000000000000110010","111111111111110101","111111111111111110","000000000000000010","111111111111010100","111111111111110100","111111111111111101","000000000000001111","111111111111010010"),
("000000000000001011","000000000000011010","111111111110110110","000000000000010110","111111111110101000","111111111111110111","000000000000011100","000000000000010011","000000000000000000","000000000000101110","111111111111101000","000000000000001010","111111111111110000","111111111111000010","000000000000000001","000000000000100000","111111111111100111","000000000000100000","000000000000010001","000000000000010000","111111111111010101","111111111111100111","000000000000010100","111111111111100010","111111111111101001","111111111111111110","111111111111110001","111111111111111100","111111111111110000","111111111111100111","000000000000000000","000000000000001000","111111111111111110","000000000000010110","111111111111110101","111111111111101000","111111111111110101","000000000000001111","111111111111110100","111111111111110011","000000000000100110","111111111111001011","111111111111110000","111111111111111100","111111111111110100","111111111111101101","000000000000011011","000000000000011100","111111111111111101","000000000000000001","000000000000011100","111111111111100110","000000000000001110","111111111111010101","000000000000000101","111111111111000111","111111111111111101","000000000000001111","000000000000000010","111111111111111111","000000000000000000","000000000000010101","000000000000010101","111111111111100010","111111111111010011","111111111111101110","111111111111100111","000000000000011111","111111111111011000","111111111111110111","000000000000011111","000000000000010100","111111111111100001","000000000000010100","000000000000010111","111111111111110110","111111111111101111","000000000000010101","111111111111111001","111111111111100000","111111111111010110","000000000000000101","111111111111100001","111111111110101111","000000000000000101","111111111111001010","111111111111001101","000000000000001100","111111111111110100","111111111111111001","000000000000011100","000000000000001011","000000000000010010","000000000000101110","111111111111000011","000000000000011111","111111111111110000","111111111111110111","111111111111111010","000000000000000110","000000000000011000","000000000000011110","111111111111110010","000000000000001100","111111111111110110","000000000000101000","111111111110110001","000000000000100111","111111111111000001","111111111111100001","111111111111100100","111111111111111100","111111111111111000","000000000000001000","111111111110011101","000000000000110110","000000000000010010","000000000000000010","111111111110111100","000000000000101010","111111111111111001","111111111111110000","111111111111110111","111111111111101011","111111111111100010","000000000000011100","111111111111110100","111111111111011111"),
("111111111111110100","000000000000010110","111111111111011010","000000000000010110","111111111110001000","111111111111110010","000000000000010111","111111111111110010","111111111111110110","000000000000110001","111111111111101001","111111111111101101","111111111110111110","111111111110101011","000000000000011010","000000000000001001","000000000000100011","000000000000010000","111111111111100110","000000000000100110","111111111111000111","111111111111111000","000000000000001100","111111111111100101","111111111111101001","000000000000001001","111111111111100000","111111111111110001","111111111111011100","111111111111001101","000000000000000110","000000000000011001","000000000000010100","111111111111111111","111111111111111110","111111111111110010","111111111111100010","111111111111110001","000000000000000010","000000000000011010","000000000000100010","111111111111101001","111111111111101110","000000000000001000","111111111111111001","000000000000000001","111111111111111111","111111111111111011","000000000000000000","000000000000000110","000000000000011000","000000000000010011","000000000000011100","111111111111001000","000000000000001111","111111111111001001","111111111111111000","000000000000010011","000000000000000000","000000000000000110","000000000000011110","000000000000111010","000000000000110110","111111111111011010","111111111110110011","111111111111100111","111111111111100110","000000000000011000","111111111111100000","111111111111111100","111111111111110101","000000000000000011","111111111110111010","000000000000000000","000000000000010101","111111111111111111","111111111111110111","000000000000110100","111111111111110101","000000000000001100","111111111111110000","000000000000001010","000000000000001001","111111111110111010","000000000000010100","111111111111111101","111111111111011100","111111111111110010","000000000000011101","111111111111111101","000000000000100011","000000000000000000","000000000000010110","000000000000010011","111111111111001100","000000000000110000","111111111111101100","111111111111111001","111111111111111110","000000000000001010","111111111111111100","000000000000000000","000000000000001101","000000000000001100","111111111110111111","000000000000010001","111111111110110010","000000000000101100","111111111111000111","111111111111101011","111111111111100011","111111111111110111","000000000000011100","000000000000001100","111111111110111001","000000000000100101","000000000000011000","000000000000000010","111111111111011000","000000000000000100","111111111111111000","111111111111101111","000000000000001010","111111111111101000","000000000000000010","000000000000001001","111111111111101011","111111111111011001"),
("111111111111011110","000000000000011110","111111111111001111","000000000000000011","111111111110010001","000000000000001110","000000000000011100","111111111111101110","000000000000000010","000000000000001100","111111111111010111","111111111111100011","111111111111001100","111111111110101010","111111111111100101","000000000000000000","000000000000001110","000000000000001100","111111111111101101","000000000000010000","111111111111001110","111111111111111100","000000000000101010","111111111111100101","111111111111101111","000000000000000100","111111111111101100","111111111111101110","111111111111110111","111111111111011111","000000000000010111","000000000000010010","000000000000000001","000000000000001001","000000000000000010","111111111111110001","111111111111011111","000000000000001100","111111111111111001","000000000000001001","000000000000011110","111111111111110111","111111111111100111","111111111111110110","000000000000001011","000000000000010001","111111111111101010","000000000000010101","000000000000000010","111111111111101110","000000000000000000","111111111111101100","111111111111111111","111111111111100101","000000000000000001","111111111111101011","000000000000000010","000000000000001000","000000000000001100","000000000000000110","000000000000101101","000000000000101110","000000000000001101","111111111111000101","111111111111000101","111111111111111110","111111111111101010","000000000000010101","111111111111100111","000000000000010011","000000000000001010","000000000000000000","111111111111000000","111111111111100110","000000000000100101","111111111111111100","111111111111100111","000000000000100111","111111111111011010","000000000000000100","111111111111110010","111111111111111011","000000000000000010","111111111111001011","000000000000000100","111111111111100101","000000000000001010","000000000000000001","000000000000001110","000000000000001011","111111111111111000","000000000000000000","000000000000011000","000000000000010000","111111111111010000","000000000000011111","111111111111111010","000000000000011100","000000000000001011","000000000000000100","111111111111111100","000000000000000000","111111111111110111","000000000000001100","111111111111011011","111111111111111101","111111111111100011","000000000000110011","111111111111100001","111111111111100010","111111111111101010","000000000000000110","000000000000011001","000000000000011101","111111111111110010","000000000000001000","000000000000000001","000000000000011101","111111111111101001","000000000000001011","111111111111101100","000000000000001111","111111111111111100","111111111111011110","111111111111110000","000000000000011111","111111111111110101","111111111111101111"),
("000000000000000111","000000000000011000","111111111111101000","000000000000001110","111111111110111110","111111111111111111","000000000000000000","111111111111110000","000000000000010000","000000000000110000","111111111111100101","111111111111101111","111111111111100110","111111111110111000","111111111111110010","000000000000000000","000000000000011011","000000000000011101","111111111111101011","000000000000011100","111111111111101001","000000000000000110","000000000000100001","111111111111011100","111111111111100001","000000000000011001","111111111111110010","111111111111111110","000000000000001001","000000000000001011","000000000000010011","000000000000011010","000000000000000110","111111111111111110","111111111111111111","111111111111110001","000000000000000000","111111111111111111","111111111111011110","111111111111111101","000000000000011110","000000000000001000","111111111111011110","000000000000000111","111111111111110000","000000000000001111","111111111111111100","000000000000001100","111111111111111100","111111111111100010","000000000000010000","000000000000000011","111111111111110110","111111111111101001","000000000000010000","111111111111100111","000000000000000000","111111111111110100","111111111111111010","000000000000000001","000000000000011101","000000000000100010","000000000000101100","111111111110101110","111111111111000110","111111111111011011","000000000000000011","000000000000010010","111111111111101111","111111111111101111","000000000000001000","000000000000010110","111111111111010110","111111111111010010","000000000000010101","111111111111101100","111111111111111001","000000000000010011","111111111111010001","000000000000001001","111111111111010010","111111111111100011","000000000000001101","111111111110111110","000000000000100101","111111111111101010","111111111111100000","000000000000001001","000000000000010000","000000000000001100","000000000000001010","111111111111111001","111111111111010011","000000000000000100","111111111111010111","000000000000100000","111111111111101000","000000000000010101","000000000000000001","111111111111011100","000000000000001100","111111111111101111","000000000000100111","000000000000010101","111111111111010011","000000000000000100","111111111111100001","000000000000001101","111111111111100100","111111111111111010","111111111111101000","000000000000000010","000000000000000101","000000000000001100","111111111111110011","000000000000101101","000000000000010101","111111111111101110","111111111111000011","111111111111100111","111111111111011101","000000000000000001","000000000000000001","111111111111011000","111111111111110001","000000000000001110","000000000000000111","111111111111111000"),
("111111111111110000","000000000000010011","000000000000010011","000000000000001000","111111111111111100","111111111111110111","000000000000001100","111111111111101001","111111111111111111","000000000000100000","111111111111010010","111111111111101011","111111111111101101","111111111110111110","000000000000001101","111111111111111010","111111111111101101","111111111111111111","111111111111100101","000000000000001110","111111111111110101","000000000000011011","111111111111111010","111111111111011000","000000000000000000","111111111111110100","111111111111011001","111111111111100111","111111111111110010","000000000000100010","000000000000010000","000000000000000010","111111111111110101","000000000000101110","000000000000000100","111111111111111110","000000000000011011","000000000000000111","111111111111010110","000000000000001010","111111111111110110","000000000000001101","111111111111101101","111111111111100100","111111111111111100","000000000000010110","111111111111101101","000000000000000011","000000000000000010","111111111111101000","000000000000100100","000000000000001010","000000000000000111","111111111111011011","000000000000000101","111111111111011000","111111111111101101","000000000000000100","111111111111111010","111111111111110000","000000000000010000","000000000001000000","000000000000001010","111111111111001000","111111111110110010","111111111111111010","000000000000011010","000000000000010111","111111111111111111","000000000000001011","000000000000010110","000000000000011111","000000000000011000","111111111111000100","000000000000000001","111111111111111011","111111111111110110","000000000000000111","111111111111010100","111111111111110100","111111111111010000","000000000000000000","111111111111101111","111111111110110111","000000000000010010","111111111111011100","000000000000000000","000000000000011001","000000000000000000","111111111111100111","111111111111111100","000000000000000010","111111111111100001","000000000000010111","111111111111110011","000000000000011000","111111111111111110","000000000000010001","000000000000000100","000000000000000000","111111111111111111","111111111111110111","000000000000010100","000000000000000001","111111111111101101","000000000000000001","111111111111111000","111111111111111011","111111111111110011","111111111111011110","111111111111110101","111111111111110001","111111111111101110","111111111111111110","111111111111110011","000000000000011101","111111111111111011","111111111111101011","111111111111110011","111111111111110101","111111111111011111","111111111111100000","111111111111111111","111111111111110100","111111111111110010","000000000000100011","000000000000000111","111111111111111001"),
("111111111111111000","000000000000010001","000000000000100101","000000000000001010","000000000000000001","000000000000001011","111111111111101101","111111111111111101","111111111111111001","111111111111101111","111111111111100001","111111111111110010","111111111111100111","111111111111001001","111111111111110111","000000000000000110","111111111111110111","000000000000001111","000000000000010110","000000000000010110","111111111111110111","111111111111110110","111111111111011110","111111111111100010","111111111111110101","000000000000001100","000000000000001100","111111111111001110","111111111111110110","000000000000000100","000000000000010100","000000000000011111","000000000000001011","000000000000101011","111111111111101110","000000000000011001","000000000000010001","000000000000000001","111111111111010101","111111111111111101","000000000000001000","000000000000010000","111111111111011101","111111111111100110","000000000000001100","000000000000000001","111111111111111000","000000000000010011","000000000000000000","111111111111101111","111111111111101100","111111111111101100","000000000000010001","111111111111111011","111111111111101101","111111111111100101","111111111111101011","111111111111101011","111111111111100110","111111111111110011","000000000000101010","000000000000101101","111111111111110001","111111111111010000","111111111110111110","000000000000010101","000000000000101000","000000000000010010","000000000000010111","000000000000000010","000000000000010100","000000000000010011","000000000000000111","111111111111001101","000000000000010101","000000000000000111","111111111111110110","000000000000000001","111111111111010001","111111111111101000","111111111111001110","000000000000001001","111111111111010111","111111111111100100","000000000000000011","111111111110111010","111111111111110100","000000000000011101","000000000000010011","111111111111011010","000000000000011100","000000000000100000","000000000000000100","000000000000001001","111111111111101011","000000000000101111","111111111111010011","000000000000000111","000000000000100100","111111111111011100","000000000000001000","000000000000001111","000000000000100010","000000000000010011","111111111111011100","111111111111110111","000000000000001111","000000000000000100","000000000000000010","111111111111010100","000000000000001000","000000000000011110","000000000000011001","000000000000011011","111111111111111110","000000000000001100","000000000000010100","111111111111011100","111111111111100010","111111111111101111","000000000000010001","111111111111100100","111111111111010011","000000000000000001","111111111111001100","000000000000110000","000000000000000000","000000000000000110"),
("111111111111111100","000000000000000111","000000000000001110","111111111111100111","000000000000010100","000000000000001000","111111111111111010","000000000000001010","111111111111010110","000000000000000000","000000000000000010","000000000000001111","000000000000001101","111111111111011100","111111111111110000","000000000000000100","111111111111110111","000000000000000101","000000000000011000","111111111111110011","111111111111101100","000000000000001010","111111111111100100","111111111111101010","111111111111111111","111111111111111111","000000000000000100","111111111111101101","111111111111100011","000000000000010000","111111111111111000","000000000000011100","000000000000000101","000000000000101001","111111111111110011","111111111111110101","000000000000010010","111111111111111100","111111111111101100","111111111111111011","111111111111110110","111111111111111100","111111111111110111","111111111111110100","000000000000001000","000000000000001000","000000000000000000","000000000000100110","000000000000011011","111111111111111001","111111111111100000","111111111111110001","000000000000000110","111111111111101010","111111111111111110","111111111111100100","111111111111110001","000000000000000011","111111111111101001","000000000000000100","000000000000000100","000000000000011101","111111111111101011","111111111111010010","111111111111100111","111111111111110110","000000000000000011","000000000000011110","000000000000000011","000000000000001000","000000000000010001","000000000000011100","000000000000010000","111111111111000111","000000000000011111","000000000000010010","000000000000010000","111111111111110010","111111111111100111","111111111111011101","111111111111110101","000000000000000110","111111111111100001","111111111111111000","111111111111111100","111111111111011000","000000000000000010","000000000000110010","000000000000000000","000000000000001100","000000000000000010","000000000000010001","111111111111100100","111111111111100011","111111111111111001","000000000000001010","111111111111011110","000000000000001110","000000000000011010","111111111111101010","111111111111111000","111111111111110011","000000000000010011","000000000000011010","111111111111010010","111111111111011111","111111111111111101","111111111111110110","111111111111110111","111111111111101100","111111111111100110","000000000000010010","000000000000000001","000000000000001001","000000000000011011","111111111111111101","000000000000010111","111111111111110010","111111111111110011","000000000000001100","000000000000100000","111111111111011011","111111111111011101","000000000000000000","111111111111110011","000000000000100011","111111111111111110","000000000000001010"),
("111111111111111010","111111111111111101","000000000000000101","111111111111110001","000000000000001010","111111111111101000","111111111111011101","111111111111110011","111111111111101110","111111111111111110","111111111111011111","000000000000000011","111111111111111010","111111111111110011","111111111111100110","111111111111100101","111111111111110011","111111111111111110","000000000000010101","000000000000000001","111111111111100000","000000000000011101","111111111111011011","111111111111001001","111111111111110101","111111111111100011","000000000000001001","111111111111101110","000000000000000110","000000000000000001","111111111111110100","000000000000010110","000000000000001100","000000000000000011","111111111111111111","000000000000011101","000000000000000001","000000000000011010","111111111111111001","000000000000011100","000000000000010000","111111111111101101","000000000000000010","111111111111101001","000000000000011011","000000000000000110","111111111111111011","111111111111110011","000000000000110101","000000000000000010","000000000000000100","111111111111111000","111111111111101010","111111111111110000","000000000000001000","111111111111100000","111111111111111000","111111111111110110","111111111111101001","000000000000001100","000000000000110111","000000000000010001","111111111111110100","111111111111011000","111111111111001010","000000000000010110","000000000000001111","111111111111110100","111111111111011011","000000000000010111","111111111111110101","000000000000010010","000000000000011100","111111111111010101","000000000000100010","000000000000001110","111111111111101101","000000000000000011","111111111111111010","111111111111101010","111111111111101110","000000000000010001","111111111111010001","111111111111101110","111111111111111101","111111111111101001","000000000000001011","000000000000010111","111111111111111000","111111111111111100","111111111111110110","000000000000000011","111111111111100000","111111111111101000","111111111111110110","111111111111110101","111111111111111001","000000000000010110","000000000000010100","000000000000010100","111111111111111110","000000000000000011","000000000000101001","000000000000000101","111111111111000011","111111111111011111","111111111111101010","111111111111111010","111111111111101010","111111111111111111","111111111111011110","000000000000000000","111111111111110010","000000000000101101","000000000000000101","111111111111111011","000000000000010010","111111111111110101","111111111111011010","000000000000010100","000000000000100000","111111111111101011","111111111111110000","111111111111100001","111111111111011111","000000000000100101","111111111111101111","000000000000011001"),
("000000000000001010","111111111111101100","000000000000001010","000000000000000000","000000000000000111","111111111111111100","000000000000000100","111111111111111110","111111111111110000","111111111111100101","111111111111011111","111111111111110101","111111111111111000","111111111111101010","000000000000000110","111111111111101100","111111111111101001","111111111111110110","000000000000001000","111111111111110110","111111111111100011","000000000000100100","111111111111110110","111111111111010111","111111111111110110","000000000000001001","000000000000011010","111111111111010011","111111111111111001","000000000000000101","111111111111111000","111111111111101110","000000000000001000","000000000000110100","111111111111111111","000000000000000010","000000000000010011","111111111111110011","111111111111110010","000000000000000111","000000000000010110","000000000000011111","000000000000000100","111111111111100111","000000000000011010","000000000000000010","000000000000000101","000000000000111011","000000000000001100","111111111111111110","111111111111011110","111111111111110001","111111111111110100","111111111111110011","111111111111111000","111111111111010101","000000000000101101","111111111111101110","111111111111101111","000000000000000000","000000000000010011","111111111111110111","111111111111110100","111111111111011100","111111111110111011","000000000000001111","000000000000001101","000000000000010010","000000000000010000","000000000000101111","111111111111110100","111111111111110110","000000000000100011","111111111111010000","000000000000110000","000000000000001000","000000000000101000","111111111111101101","111111111111111101","111111111111111000","000000000000010011","000000000000010010","111111111111111101","111111111111011110","111111111111111000","111111111111101000","000000000000010111","000000000000000010","000000000000001110","000000000000000000","111111111111101011","000000000000000111","000000000000000101","111111111111100100","000000000000000001","000000000000001110","111111111111101111","000000000000011100","000000000000011101","000000000000011011","000000000000010001","000000000000101010","000000000000000010","111111111111110101","111111111111111010","111111111111110101","111111111111100101","111111111111011111","111111111111101010","000000000000010001","000000000000001001","111111111111101111","000000000000000001","000000000000000010","000000000000010110","111111111111110001","000000000000001001","000000000000001001","111111111111101101","111111111111101100","000000000000001010","000000000000001011","111111111111101101","111111111111011010","000000000000000001","000000000000101000","000000000000000011","000000000000001000"),
("000000000000001110","111111111111100001","111111111111111111","111111111111100110","000000000000001010","000000000000001101","000000000000001011","000000000000011010","111111111111110110","111111111111100100","000000000000001001","000000000000000000","000000000000000111","111111111111110111","111111111111110111","111111111111110101","111111111111011101","000000000000001111","000000000000100101","111111111111111010","111111111111100011","000000000000000101","111111111111110001","111111111111110101","000000000000000110","111111111111111111","000000000000100110","111111111111100111","000000000000000100","000000000000000100","000000000000000110","111111111111100110","000000000000000110","111111111111111111","000000000000101000","111111111111111100","000000000000011110","111111111111101010","111111111111110011","111111111111011011","111111111111110011","000000000000011100","000000000000000010","111111111111111100","000000000000010111","111111111111110110","000000000000001001","000000000000110100","111111111111110111","000000000000000101","111111111111110010","000000000000000000","000000000000001100","111111111111011110","000000000000000000","111111111111111011","000000000000001010","111111111111101111","000000000000000001","111111111111111011","111111111111111111","111111111111110111","111111111111110001","000000000000010011","111111111111010111","000000000000000101","000000000000000011","000000000000011111","000000000000011011","000000000000001100","000000000000010000","111111111111011111","000000000000100111","111111111111111011","000000000000010000","111111111111110010","000000000000011101","111111111111110100","111111111111111000","111111111111111000","000000000000100011","111111111111111010","111111111111111011","111111111111110110","111111111111110011","000000000000000101","111111111111101010","111111111111101000","000000000000100110","111111111111101110","000000000000000010","111111111111110110","000000000000001000","111111111111111111","000000000000000011","000000000000100000","111111111111011100","000000000000000011","000000000000010110","000000000000001000","000000000000001001","000000000000110001","000000000000001101","000000000000010011","000000000000010000","000000000000010000","111111111111111011","111111111111011101","111111111111010101","000000000000000010","111111111111100001","000000000000000000","000000000000001001","111111111111101100","000000000000100010","000000000000000010","111111111111110111","000000000000000000","111111111111111110","111111111111110100","111111111111111011","000000000000001011","111111111111110100","000000000000011111","111111111111101101","111111111111111101","000000000000100111","111111111111110000"),
("111111111111111111","111111111111101111","111111111111100111","111111111111100111","000000000000011011","000000000000010100","000000000000010101","000000000000001010","000000000000001010","000000000000000100","111111111111101000","000000000000001111","000000000000000110","111111111111001011","111111111111110110","111111111111111100","000000000000001101","000000000000000110","000000000000001010","111111111111101011","111111111111010010","000000000000011100","111111111111110101","000000000000010011","000000000000000111","000000000000011011","000000000000001010","111111111111101111","000000000000101100","000000000000000010","000000000000000011","111111111111111001","000000000000000001","000000000000100101","000000000000010000","000000000000010101","000000000000000000","111111111111111100","000000000000000110","111111111111110100","000000000000000101","000000000000011101","111111111111111010","000000000000000100","000000000000000111","000000000000010010","000000000000000001","000000000000111101","000000000000010011","000000000000000010","111111111111101011","111111111111101111","000000000000001000","111111111111110010","111111111111100001","111111111111101000","000000000000011000","111111111111110010","111111111111111100","000000000000000100","000000000000001010","111111111111100101","111111111111010111","111111111111111100","111111111111101101","000000000000001001","000000000000000000","000000000000101011","111111111111110010","000000000000001001","000000000000010001","111111111111011101","000000000000110101","111111111111110101","000000000000010001","111111111111101100","000000000000001010","111111111111011101","000000000000010100","000000000000001110","000000000000010110","000000000000001010","000000000000000001","111111111111100000","111111111111111001","111111111111110110","111111111111100011","111111111111111100","000000000000011100","000000000000001101","000000000000010010","000000000000100001","111111111111101001","000000000000000001","111111111111111000","111111111111111001","111111111111110001","000000000000010100","000000000000011001","000000000000000001","000000000000011110","000000000000101101","000000000000101100","000000000000000011","111111111111101100","000000000000100010","000000000000010000","111111111111110100","111111111111011111","111111111111110110","111111111111110010","111111111111111101","000000000000001100","111111111111101011","000000000000001011","111111111111111111","000000000000010011","000000000000000010","000000000000000001","111111111111100000","000000000000001110","111111111111110100","111111111111101001","000000000000011101","000000000000000000","000000000000000000","111111111111111100","000000000000000101"),
("111111111111111110","111111111111111001","111111111111111100","000000000000000011","000000000000001001","000000000000010010","000000000000010010","000000000000001111","111111111111111100","111111111111110100","111111111111111010","111111111111110011","000000000000001110","111111111111011001","000000000000010011","000000000000000101","000000000000010110","111111111111101001","000000000000001000","111111111111011010","111111111111101010","111111111111110110","000000000000001010","000000000000001010","000000000000001010","000000000000001010","111111111111011010","111111111111111110","000000000000100101","000000000000000101","111111111111111110","111111111111101000","000000000000001101","000000000000011101","111111111111111111","000000000000000010","111111111111101110","111111111111101000","111111111111111100","111111111111111000","000000000000000110","000000000000011111","111111111111111111","000000000000010101","000000000000001101","000000000000010101","111111111111101111","000000000000001101","000000000000000010","000000000000001111","111111111111100001","000000000000000000","000000000000011110","111111111111111111","000000000000000011","111111111111101100","111111111111101000","111111111111011011","000000000000010011","111111111111110000","000000000000000100","111111111111101101","111111111111011011","111111111111110000","111111111111101101","111111111111111010","111111111111111100","000000000000010001","111111111111111110","111111111111100010","000000000000000011","111111111111110011","111111111111111111","111111111111110110","000000000000001001","000000000000001011","000000000000000001","000000000000000000","111111111111111101","000000000000001010","000000000000001000","000000000000000000","111111111111111100","111111111111011011","000000000000000110","111111111111111100","000000000000000101","111111111111101101","000000000000100001","111111111111111010","111111111111110011","000000000000000101","111111111111101101","111111111111111101","111111111111100110","000000000000101100","000000000000001000","000000000000001000","111111111111110111","111111111111100011","000000000000010110","111111111111111001","000000000000110000","111111111111100110","111111111111100111","000000000000010000","111111111111111110","111111111111101111","111111111111100011","000000000000000110","111111111111111001","111111111111111100","000000000000011001","111111111111110000","111111111111111011","000000000000010110","000000000000010110","000000000000001101","111111111111110111","111111111111111001","111111111111110010","111111111111111000","000000000000010100","000000000000000111","111111111111110110","000000000000010000","000000000000001010","111111111111110001"),
("111111111111101101","000000000000001111","111111111111101000","000000000000001010","111111111111101100","111111111111111000","000000000000000010","000000000000001000","000000000000000010","111111111111111110","000000000000011001","111111111111111000","000000000000011110","111111111111111000","111111111111111010","000000000000010110","111111111111100111","000000000000100001","000000000000001111","111111111111111011","111111111111111100","000000000000011110","000000000000000000","000000000000001111","000000000000010011","111111111111101001","111111111111111011","000000000000010000","111111111111111101","000000000000000110","000000000000010010","000000000000001100","000000000000011011","000000000000001000","111111111111111110","000000000000001100","000000000000010110","000000000000001011","000000000000000100","111111111111101100","000000000000001001","111111111111110011","000000000000010000","111111111111101010","000000000000000010","111111111111110011","111111111111111101","111111111111110111","000000000000000100","111111111111110001","111111111111111010","000000000000000111","000000000000001000","000000000000010101","111111111111111110","111111111111111110","000000000000000010","000000000000010000","111111111111111111","111111111111110001","000000000000011001","000000000000000010","111111111111100010","111111111111101100","111111111111110000","000000000000000000","111111111111111011","111111111111101011","000000000000010000","000000000000010000","111111111111100010","000000000000011100","111111111111101101","000000000000001101","111111111111111011","000000000000000000","000000000000010010","000000000000011110","000000000000010010","111111111111111001","000000000000000110","000000000000011101","111111111111111011","111111111111110001","000000000000010101","111111111111111100","111111111111111100","000000000000011101","111111111111111011","000000000000000011","111111111111101011","000000000000010010","111111111111110001","111111111111011111","000000000000001101","111111111111110100","000000000000001101","000000000000000101","000000000000001010","000000000000000001","000000000000001011","111111111111110110","000000000000001000","111111111111111110","000000000000011010","000000000000000111","000000000000000100","000000000000010110","111111111111101101","000000000000001011","000000000000000010","000000000000000000","000000000000000000","111111111111101011","111111111111111101","111111111111101000","000000000000000100","000000000000010001","000000000000000000","111111111111110101","000000000000000110","000000000000011100","000000000000010000","000000000000010111","000000000000001101","111111111111011111","000000000000100110","111111111111110010"),
("000000000000011100","000000000000001100","000000000000010011","111111111111111010","000000000000001111","000000000000000011","111111111111110100","111111111111110101","111111111111100110","111111111111011010","111111111111110011","000000000000010000","000000000000001001","000000000000001111","000000000000010000","111111111111111101","000000000000010001","000000000000000111","111111111111111001","000000000000010110","000000000000010001","111111111111111100","111111111111011001","111111111111100110","000000000000010110","111111111111101010","111111111111101011","111111111111111000","000000000000100100","000000000000001111","111111111111111011","111111111111111001","000000000000100010","111111111111110101","111111111111110110","111111111111100100","000000000000010000","000000000000001001","111111111111111010","111111111111111010","000000000000100001","000000000000011011","000000000000001111","111111111111101100","000000000000011001","111111111111110000","000000000000001000","000000000000010010","000000000000000111","000000000000010010","111111111111111100","000000000000001100","111111111111111111","000000000000010100","111111111111101011","111111111111110010","000000000000010011","000000000000000011","000000000000000111","111111111111101110","000000000000001111","111111111111111010","111111111111111110","000000000000000011","111111111111111000","000000000000001110","000000000000010000","111111111111111010","111111111111111000","111111111111111010","111111111111111011","000000000000001011","000000000000100110","111111111111111100","000000000000011000","000000000000000001","000000000000000001","000000000000000100","000000000000010110","111111111111111010","111111111111110101","000000000000000100","000000000000001111","111111111111100110","000000000000000111","000000000000011000","000000000000000000","111111111111111111","111111111111110101","111111111111110010","000000000000000011","000000000000010001","111111111111101110","111111111111100010","111111111111111110","111111111111111010","000000000000000100","111111111111111001","000000000000000000","111111111111101110","000000000000001010","111111111111111101","111111111111101111","111111111111101000","000000000000001100","111111111111101110","000000000000000000","111111111111111001","111111111111100010","000000000000010011","111111111111110001","000000000000011111","000000000000001000","111111111111110110","111111111111100001","000000000000000110","111111111111111100","111111111111111101","111111111111101001","111111111111111100","000000000000001000","000000000000010110","111111111111110011","000000000000010001","000000000000000111","111111111111101011","000000000000010001","000000000000000001"),
("111111111111110000","000000000000001110","000000000000001011","000000000000000110","000000000000000000","111111111111110010","111111111111110001","000000000000000110","111111111111111100","111111111111111001","000000000000010011","111111111111110111","000000000000001011","000000000000001001","111111111111110101","000000000000001101","000000000000001011","111111111111110111","111111111111101111","000000000000001101","111111111111111000","000000000000000010","111111111111111000","000000000000000110","000000000000000111","000000000000001000","000000000000000111","000000000000001100","111111111111110101","000000000000001010","111111111111110010","000000000000001000","000000000000001000","000000000000000010","111111111111111111","000000000000010011","111111111111111001","000000000000010011","000000000000001100","000000000000001010","111111111111111111","000000000000000010","000000000000001001","111111111111110011","111111111111110001","000000000000010001","111111111111110000","000000000000010100","111111111111110000","000000000000000010","111111111111111100","111111111111101101","000000000000001000","000000000000001111","000000000000001100","000000000000010001","000000000000000111","000000000000001110","000000000000001011","111111111111110010","000000000000010010","111111111111111110","111111111111111011","111111111111111110","000000000000010001","000000000000000100","000000000000001101","000000000000000110","000000000000000011","000000000000000100","111111111111111110","111111111111110010","000000000000000011","111111111111110100","111111111111110010","000000000000001000","000000000000001101","000000000000001110","000000000000010000","000000000000000011","111111111111101111","111111111111110110","111111111111111010","111111111111110100","111111111111111101","111111111111110000","000000000000010000","000000000000001010","000000000000001100","000000000000000000","000000000000010100","000000000000000000","111111111111111001","111111111111110000","000000000000010010","111111111111110111","000000000000000000","111111111111111100","000000000000000110","000000000000000110","111111111111111011","000000000000001101","000000000000000011","111111111111111000","000000000000010001","111111111111111011","000000000000010000","000000000000000000","111111111111111111","111111111111111111","111111111111110001","111111111111111101","111111111111111011","000000000000010001","000000000000000000","000000000000001100","000000000000001001","111111111111111001","111111111111110101","111111111111111011","000000000000001001","111111111111101101","000000000000000111","000000000000001001","111111111111110111","000000000000000100","111111111111110010","000000000000010010"),
("111111111111110101","111111111111111010","000000000000001111","111111111111111101","111111111111101111","000000000000000110","000000000000000000","111111111111110110","111111111111110100","000000000000000101","111111111111101111","111111111111111111","000000000000001111","000000000000001000","000000000000000101","000000000000001010","000000000000001100","000000000000000111","000000000000001111","000000000000001000","111111111111110111","111111111111110000","000000000000010000","000000000000000111","000000000000000000","111111111111111101","111111111111110010","000000000000000101","111111111111110111","000000000000000000","000000000000001010","111111111111101100","111111111111111111","000000000000001011","111111111111101101","000000000000001000","000000000000000000","000000000000000000","000000000000001011","111111111111110110","111111111111111110","000000000000010010","000000000000001000","000000000000000001","000000000000010010","000000000000000110","111111111111110101","111111111111111001","000000000000000000","111111111111110100","111111111111110001","000000000000010100","111111111111111101","111111111111111111","111111111111111111","111111111111111101","000000000000001110","111111111111110110","000000000000000110","111111111111110010","111111111111111100","111111111111110011","000000000000000000","111111111111111111","000000000000010011","111111111111111001","111111111111101111","000000000000010001","000000000000000000","111111111111110001","000000000000010000","111111111111111110","000000000000000000","111111111111110110","000000000000000100","000000000000000000","111111111111110001","000000000000001110","111111111111111001","111111111111101100","000000000000001000","000000000000000010","000000000000001011","111111111111111000","111111111111111110","111111111111110010","111111111111111111","000000000000010100","111111111111110001","111111111111111110","000000000000000110","000000000000000011","111111111111101101","111111111111111110","111111111111110110","111111111111101111","000000000000000011","000000000000000100","111111111111110000","111111111111101100","111111111111111110","111111111111110101","000000000000001010","000000000000001011","000000000000000000","000000000000001101","000000000000001000","000000000000000000","111111111111111010","000000000000001110","000000000000000011","111111111111110000","111111111111101101","000000000000001111","000000000000001101","111111111111111010","111111111111111110","000000000000001100","111111111111110010","111111111111111100","111111111111110110","000000000000010001","000000000000001000","111111111111111101","111111111111101101","111111111111110110","000000000000001001","111111111111110110"),
("111111111111101101","111111111111110111","111111111111110110","000000000000001000","111111111111111101","000000000000000011","111111111111110101","000000000000001010","000000000000001101","000000000000001010","000000000000001011","000000000000000101","111111111111111010","000000000000000111","000000000000000110","000000000000000010","111111111111101110","000000000000000011","000000000000000101","000000000000000010","111111111111110011","000000000000010001","000000000000000011","111111111111111111","111111111111111001","111111111111110000","000000000000000011","111111111111111111","000000000000010010","000000000000000011","111111111111111101","000000000000010001","000000000000001000","000000000000000111","000000000000000111","000000000000001000","111111111111110000","111111111111111110","000000000000001010","000000000000000110","111111111111111100","000000000000001111","000000000000000101","000000000000010000","000000000000000100","111111111111111011","111111111111110110","111111111111110010","111111111111111110","111111111111111101","000000000000000111","111111111111111111","111111111111110111","111111111111101110","000000000000001101","000000000000000011","000000000000000000","000000000000001010","111111111111110110","111111111111111100","000000000000001101","000000000000000100","111111111111101110","000000000000000011","111111111111111001","000000000000000111","000000000000000011","111111111111110010","000000000000001000","000000000000000010","000000000000000111","000000000000001001","111111111111110011","111111111111111011","111111111111110111","000000000000000111","111111111111110110","000000000000010100","000000000000010000","000000000000010011","000000000000001111","111111111111111000","111111111111110100","000000000000000000","000000000000010010","000000000000001110","111111111111111000","000000000000010010","000000000000001000","000000000000000100","111111111111111001","000000000000010101","111111111111101110","000000000000000001","111111111111110001","000000000000000000","000000000000000000","111111111111111000","000000000000000110","000000000000000001","111111111111111000","111111111111111111","000000000000000101","000000000000000010","000000000000000111","000000000000000101","000000000000010011","111111111111111100","000000000000001111","111111111111101100","000000000000010100","000000000000010000","111111111111111110","111111111111110010","111111111111110101","111111111111111111","000000000000001011","111111111111110100","111111111111101101","111111111111110010","111111111111101011","111111111111101111","000000000000000011","000000000000000110","111111111111110001","000000000000000000","000000000000000000","111111111111110101"),
("111111111111011100","111111111111111001","111111111111110000","000000000000010011","000000000000100101","111111111111101101","111111111111110011","111111111111110000","000000000000001001","111111111111111001","000000000000101110","000000000000011000","000000000000000111","000000000000000101","111111111111110011","111111111111100100","111111111111110011","000000000000001110","000000000000000101","000000000000001000","000000000000011000","111111111111100010","111111111111111010","000000000000001001","111111111111111100","000000000000000010","000000000000001000","000000000000000101","000000000000000010","000000000000000111","000000000000000000","111111111111100101","111111111111101001","000000000000000010","000000000000000110","000000000000010000","111111111111011101","000000000000011100","111111111111110000","000000000000000000","000000000000001000","000000000000000111","111111111111101010","000000000000100111","111111111111110111","000000000000110000","111111111111111011","000000000000000000","111111111111010101","111111111111101010","000000000000001110","111111111111100100","000000000000000000","000000000000011000","000000000000011101","000000000000011100","111111111111100110","000000000000000000","111111111111111000","000000000000001010","111111111111101111","000000000000010100","000000000000001110","000000000000000000","000000000000010110","111111111111100101","111111111111111000","111111111111110110","000000000000000011","000000000000000011","000000000000000100","000000000000001100","111111111111011010","000000000000010111","000000000000000111","111111111111110101","111111111111101010","000000000000000011","000000000000001100","111111111111101111","000000000000100100","111111111111100100","000000000000011001","000000000000010010","000000000000101100","111111111111110011","111111111111111101","111111111111110100","111111111111010111","000000000000100010","000000000000100110","111111111111111101","000000000000000000","000000000000100010","000000000000000110","111111111111110111","000000000000001110","111111111111101101","111111111111110110","000000000000000000","111111111111100111","000000000000001001","111111111111101111","000000000000001111","000000000000011110","111111111111011000","000000000000100010","111111111111110111","000000000000001111","000000000000000111","000000000000001100","000000000000000011","111111111111111011","111111111111111110","000000000000101011","111111111111100010","111111111111010111","000000000000100110","000000000000001100","000000000000011000","111111111111111111","000000000000001010","111111111111101101","000000000000010010","111111111111111111","111111111111010101","111111111111111010","000000000000000111"),
("111111111111101101","000000000000001101","000000000000000011","000000000000001001","000000000000001110","111111111111010101","000000000000010000","000000000000000100","000000000000000100","000000000000011010","111111111111101101","000000000000000001","000000000000000101","000000000000010000","000000000000000101","111111111111011101","111111111111100100","111111111111100101","111111111111111111","000000000000000000","000000000000001000","000000000000000110","111111111111110101","111111111111111011","111111111111111011","000000000000000111","111111111111110000","000000000000000001","000000000000001110","000000000000000111","000000000000000100","000000000000000000","000000000000000000","000000000000010011","111111111111110101","000000000000100100","000000000000000000","000000000000010101","111111111111111001","000000000000000010","000000000000000000","000000000000000011","000000000000011101","111111111111101010","111111111111101011","000000000000100100","000000000000000110","111111111111100011","000000000000000001","111111111111111101","000000000000000000","111111111111101111","000000000000011101","000000000000100111","000000000000110011","111111111111111011","111111111111101011","000000000000000111","111111111111111000","111111111111111110","111111111111111111","000000000000101100","111111111111101111","111111111111100001","000000000000101001","111111111111110100","000000000000101001","000000000000010100","000000000000001100","000000000000001000","000000000000010101","000000000000101011","111111111111110100","000000000000001011","000000000000011110","000000000000010000","111111111111101000","000000000000011011","111111111111100010","111111111111111010","111111111111111010","111111111111111111","111111111111101000","000000000000011010","000000000000010010","111111111111100110","111111111111111100","000000000000101100","000000000000001001","000000000000100101","111111111111110010","000000000000100101","000000000000000000","000000000000100011","111111111111011100","111111111111111001","000000000000001110","000000000000010000","000000000000001001","111111111111100111","111111111111111010","111111111111101101","111111111111110110","111111111111111000","000000000000010101","111111111111110101","111111111111111101","111111111111111111","000000000000010000","111111111111100010","111111111111100111","111111111111111111","000000000000010100","000000000000000000","000000000000000110","000000000000000000","000000000000000010","000000000000010010","000000000000000000","000000000000011000","000000000000001011","111111111111101011","111111111111111111","111111111111100011","111111111111010111","000000000000010010","111111111111011010","000000000000010111"),
("111111111111100101","000000000000001110","111111111111111011","111111111111111000","111111111111110010","000000000000011100","111111111111110110","000000000000001011","111111111111110000","000000000000011100","000000000000000010","000000000000000010","000000000000001101","111111111111111110","000000000000100110","111111111111110101","000000000000001110","111111111111011011","111111111111100110","111111111111101001","111111111111110110","111111111111101001","000000000000000100","000000000000000100","000000000000000111","000000000000001001","111111111111110100","000000000000001100","000000000000100000","000000000000000100","111111111111110000","000000000000011011","111111111111110100","111111111111100110","111111111111111100","000000000000011110","000000000000000000","111111111111110101","000000000000001110","111111111111101011","000000000000010010","111111111111100001","000000000000000111","111111111111110011","111111111111111011","000000000000011011","000000000000001000","111111111111101110","111111111111110001","000000000000011110","000000000000001111","111111111111101110","111111111111101101","000000000000010010","111111111111110110","111111111111111010","111111111111100101","111111111111111010","000000000000000001","000000000000001100","000000000000010101","111111111111111110","111111111111111001","111111111111111011","111111111111111100","111111111111100011","000000000000100011","000000000000001000","000000000000000110","111111111111100100","000000000000001100","000000000000000010","000000000000110000","000000000000100011","000000000000011011","111111111111111101","111111111111111000","111111111111111101","000000000000001010","111111111111111101","000000000000000001","111111111111110111","000000000000100011","000000000000011001","000000000000001110","111111111111111000","111111111111101010","000000000000100000","000000000000101000","000000000000001110","000000000000010011","000000000000011111","111111111111111111","000000000000000010","111111111111101100","000000000000001010","000000000000001001","000000000000001100","111111111111111110","000000000000000011","000000000000010111","000000000000000000","000000000000000001","111111111111111010","000000000000000101","111111111111110000","111111111111110011","000000000000100010","000000000000100010","000000000000011000","111111111111111001","111111111111111101","000000000000010101","000000000000000111","111111111111111000","000000000000010000","000000000000100011","000000000000010000","000000000000001101","111111111111110111","111111111111100111","000000000000000011","111111111111101000","000000000000101001","000000000000000000","111111111111100011","111111111111101010","000000000000001110"),
("111111111111101101","111111111111101011","111111111111100101","000000000000001000","000000000000110100","000000000000010101","111111111111110000","000000000000001111","111111111111111010","000000000000010010","111111111111111011","111111111111001101","000000000000010011","111111111111100100","000000000000011010","000000000000010101","000000000000100110","111111111111111111","000000000000100011","111111111111111111","111111111111010111","111111111111110010","111111111111110000","111111111111010001","111111111111101111","000000000000110101","000000000000000011","111111111111110110","000000000000110001","000000000000001000","000000000000000111","000000000000011111","000000000000000101","111111111111011011","111111111111110110","000000000000010111","111111111111011110","000000000000001001","000000000000000010","111111111111110100","111111111111110010","111111111111011010","000000000000100110","000000000000011100","111111111111110101","000000000000001101","000000000000011010","111111111111101011","111111111111111111","000000000000011000","111111111111111101","111111111111100100","111111111111010101","111111111111111101","111111111111110101","111111111111110101","111111111111011001","000000000000010001","111111111111110101","111111111111101100","000000000000001101","111111111111110001","000000000000000010","111111111111110010","111111111111101000","111111111111101110","000000000000010111","000000000000011100","111111111111011100","111111111111100101","000000000000010001","000000000000001111","000000000000100110","000000000000001010","000000000000100100","000000000000011001","111111111111111111","000000000000010110","000000000000001101","000000000000010101","111111111111110011","111111111111111000","000000000000100001","111111111111011111","000000000000010011","111111111111110101","111111111111100111","000000000000010101","111111111111111110","000000000000011011","000000000000000010","000000000000000001","111111111111110101","000000000000000011","111111111111101001","000000000000101111","000000000000011001","111111111111100100","111111111111110001","000000000000001000","000000000000000100","111111111111100001","000000000000010010","111111111111111110","111111111111101001","000000000000010001","000000000000000000","000000000000000010","111111111111101110","111111111111110111","111111111111100101","111111111111101011","111111111111111101","000000000000010001","111111111111011100","000000000000010010","000000000000101000","000000000000000111","111111111111110000","000000000000000101","111111111111100000","111111111111101111","000000000000010000","000000000000000010","000000000000001011","111111111111110001","000000000000001010","111111111111111011"),
("111111111111101010","111111111111110001","111111111111000010","111111111111111000","000000000000001000","000000000000110001","000000000000011101","000000000000001001","000000000000010001","111111111111110111","000000000000000001","111111111111101101","000000000000100010","111111111111111101","000000000000101100","000000000000001011","000000000000010000","000000000000000000","000000000000100100","000000000000001111","111111111111000100","111111111111001011","111111111111100111","111111111111100110","111111111111110101","000000000000110011","000000000000010010","000000000000100001","000000000000110000","111111111111110011","000000000000010000","000000000000000011","000000000000000011","111111111111010111","000000000000000011","000000000000011001","111111111111110111","000000000000000110","111111111111111110","111111111111111101","000000000000001010","111111111111101001","000000000000100110","000000000000000111","000000000000000101","111111111111111000","000000000000011101","000000000000000111","111111111111011011","000000000000001001","000000000000100010","111111111111101000","111111111111100100","111111111111111001","000000000000000000","111111111111110000","111111111111100000","000000000000000010","111111111111100101","000000000000010001","111111111111110100","000000000000010001","000000000000011101","000000000000000000","000000000000010000","111111111111100110","000000000000010110","000000000000010000","111111111111111100","111111111111011011","000000000000110001","000000000000100010","000000000000000010","111111111111111001","000000000000001111","000000000000100010","000000000000001100","000000000000000100","000000000000000011","000000000000000000","111111111111100111","000000000000001010","000000000000111011","111111111111010101","111111111111111010","111111111111101011","111111111111111000","000000000000010111","111111111111101110","000000000000001001","111111111111110010","111111111111111100","111111111111110111","000000000000000000","111111111111100101","000000000000010001","000000000000010001","000000000000010011","111111111111110000","111111111111011001","000000000000001101","000000000000000000","000000000000000101","000000000000011101","111111111111011110","000000000000001101","111111111111011101","000000000000000000","111111111111111011","111111111111101110","111111111111011101","000000000000001100","111111111111110110","111111111111111101","111111111111011000","000000000000100001","000000000000001111","000000000000000101","111111111111101010","000000000000001000","000000000000010000","111111111111100001","111111111111100001","000000000000010110","000000000000101100","111111111111110010","000000000000010001","111111111111101000"),
("111111111111010010","000000000000000101","111111111111000010","111111111111101111","000000000000010111","000000000000100000","111111111111110110","000000000000010000","111111111111111111","111111111111100110","111111111111111111","111111111111101001","111111111111111010","111111111111111000","000000000000011000","000000000000010000","000000000000000110","000000000000010001","000000000000011111","111111111111111111","111111111110111000","111111111111100011","111111111111110100","111111111111110110","111111111111110101","000000000000000001","000000000000001111","000000000000010100","000000000000000101","111111111111110001","000000000000000101","000000000000001100","000000000000001001","111111111111100001","000000000000000101","000000000000001011","111111111111111111","000000000000010000","111111111111100010","000000000000000101","111111111111111101","111111111111001100","000000000000010100","000000000000011110","000000000000001110","111111111111110100","000000000000100000","000000000000011100","000000000000000101","111111111111111101","111111111111111001","000000000000010010","111111111111111000","000000000000001101","000000000000000000","000000000000000010","111111111111011011","000000000000000011","111111111111110001","111111111111111111","111111111111110000","000000000000011010","000000000000001010","000000000000000100","111111111111101100","111111111111110111","111111111111110100","000000000000001101","111111111111110000","111111111111110111","000000000000011110","000000000000010010","000000000000001010","000000000000001110","000000000000100100","000000000000010101","111111111111101111","000000000000010111","111111111111111010","000000000000011001","000000000000000100","000000000000000011","000000000000000101","111111111111101001","000000000000001100","111111111111011110","000000000000000001","000000000000010010","111111111111101101","111111111111111010","111111111111110000","111111111111110111","000000000000000111","111111111111111110","111111111111001101","111111111111111001","111111111111110100","111111111111101111","111111111111010011","000000000000000010","000000000000010100","000000000000011000","000000000000010011","000000000000000010","111111111111101010","000000000000000010","111111111111000111","000000000000001100","111111111111100101","000000000000000101","111111111111100001","000000000000001000","000000000000011011","000000000000010110","111111111111011110","000000000000010001","000000000000011001","000000000000010001","111111111111110001","000000000000011101","000000000000001110","111111111111101111","111111111111100110","111111111111100100","000000000000010000","111111111111111010","111111111111110100","111111111111111110"),
("111111111111100000","000000000000010110","111111111111010111","000000000000010010","000000000000100111","000000000000101011","111111111111101111","000000000000001010","000000000000011011","111111111111110110","111111111111110110","111111111111100011","000000000000001011","111111111111001110","000000000000011111","000000000000001111","111111111111111101","000000000000001111","000000000000001000","000000000000010111","111111111111000000","111111111111001101","111111111111111000","111111111111110000","111111111111000111","000000000000001100","000000000000001010","000000000000100111","000000000000001101","111111111111001111","111111111111011100","000000000000010000","111111111111111100","111111111111011010","111111111111110111","000000000000011000","111111111111111111","000000000000011101","111111111111110010","111111111111111110","111111111111110101","111111111111001001","000000000000010101","000000000000100100","111111111111111101","111111111111101111","000000000000100011","000000000000010110","111111111111110001","111111111111101100","000000000000011001","111111111111111101","111111111111100001","111111111111110011","000000000000000001","111111111111011011","111111111111100101","111111111111111100","111111111111110000","111111111111111110","000000000000000000","000000000000011110","111111111111111100","111111111111111110","111111111111110100","111111111111011110","111111111111010100","000000000000101010","111111111111000101","111111111111101010","000000000000110001","000000000000100000","111111111111101001","000000000000010010","000000000000001101","111111111111111101","111111111111100110","000000000000011000","111111111111110000","000000000000010111","111111111111111011","000000000000000100","000000000000011100","111111111111100011","000000000000101011","111111111111010110","000000000000000000","000000000000010111","111111111111111011","000000000000000010","111111111111011000","000000000000001100","000000000000010001","000000000000001011","111111111111100010","111111111111110011","111111111111111111","111111111111111110","111111111111011110","111111111111110110","111111111111110000","000000000000010110","111111111111111111","000000000000001010","111111111111001111","000000000000011000","111111111111101010","000000000000010001","111111111111100011","111111111111111011","111111111111100101","111111111111110010","000000000000001001","111111111111111111","111111111111011000","000000000000001110","000000000000100001","000000000000010000","111111111111100001","000000000000011011","111111111111100101","111111111111101110","111111111111111110","000000000000000010","111111111111110001","111111111111010110","000000000000000001","111111111111110010"),
("111111111111100001","000000000000000011","111111111111000000","000000000000100001","000000000000000110","000000000000010010","111111111111110111","000000000000101010","000000000000000010","000000000000000101","000000000000000110","000000000000100010","111111111111100101","111111111111011110","000000000000001010","000000000000010110","000000000000010101","000000000000001111","000000000000100010","000000000000100011","111111111110101000","111111111111011110","111111111111111101","111111111111100010","111111111111011011","000000000000010100","000000000000000011","000000000000000000","000000000000000101","111111111111100100","111111111111111001","111111111111110111","000000000000011010","111111111111100011","111111111111111111","000000000000001010","111111111111111011","000000000000000001","111111111111110111","000000000000001001","000000000000010110","111111111111111010","111111111111111111","000000000000000110","000000000000011011","111111111111011110","000000000000101110","000000000000010011","111111111111111101","111111111111111000","000000000000101001","000000000000001011","111111111111100001","111111111111100111","000000000000010000","111111111111001011","111111111111111001","000000000000000101","111111111111110111","000000000000000110","111111111111111111","000000000000011110","000000000000100101","111111111111111000","111111111111010110","111111111111110000","111111111111001000","000000000000001010","111111111110111001","111111111111011111","000000000000011111","000000000000011110","000000000000001110","000000000000001110","000000000000000101","111111111111101011","000000000000001100","000000000000101000","111111111111101010","000000000000011011","111111111111101001","000000000000001001","000000000000010000","111111111111001011","000000000000101111","111111111111101111","000000000000000101","000000000000010100","111111111111111111","000000000000000111","111111111111101010","000000000000011001","000000000000101101","111111111111111110","111111111111100100","111111111111011000","000000000000001001","111111111111101111","111111111111001100","111111111111100101","000000000000000010","000000000000000000","000000000000000111","000000000000100010","111111111111101001","000000000000011001","111111111111010110","000000000000000101","111111111111110000","000000000000001110","111111111111101000","000000000000000001","000000000000100001","111111111111101100","111111111111011000","000000000000010001","000000000000011100","000000000000001101","111111111111010111","000000000000011001","000000000000000010","111111111111011110","111111111111110100","000000000000010000","000000000000011000","111111111111100010","111111111111101001","111111111111101000"),
("111111111111100000","000000000000100001","111111111111000111","111111111111111101","111111111111111110","000000000000011110","111111111111111110","000000000000011110","000000000000010001","000000000000001110","000000000000010010","000000000000010100","111111111111111001","111111111111000011","111111111111111100","000000000000011000","000000000000000110","111111111111111101","111111111111110011","000000000000001110","111111111111001010","111111111111111001","111111111111110101","111111111111011010","111111111111101011","000000000000001111","111111111111110011","111111111111110110","000000000000000000","111111111111010011","111111111111111100","000000000000000000","000000000000000110","111111111111110101","111111111111110000","000000000000011000","111111111111111110","000000000000100101","000000000000001011","111111111111110110","111111111111111111","000000000000000000","000000000000001100","111111111111111100","000000000000101111","111111111111011101","000000000000011100","000000000000011010","111111111111110001","000000000000000110","000000000000001000","000000000000011100","111111111111101010","111111111111111010","000000000000001111","111111111111000111","111111111111110000","111111111111111101","111111111111110101","111111111111111110","000000000000000010","000000000000011100","000000000000011000","111111111111101011","111111111111010101","111111111111101000","111111111110101100","000000000000011111","111111111110111000","111111111111001111","000000000000101111","000000000000100000","111111111111111110","111111111111111101","000000000000010111","000000000000000001","111111111111101110","000000000000010011","111111111111100101","000000000000001101","111111111111101010","000000000000000100","000000000000101110","111111111111010100","000000000000010111","111111111111011100","000000000000000001","000000000000011001","000000000000011010","000000000000001001","111111111111101111","000000000000011000","000000000000100001","111111111111111111","111111111111011000","111111111111110010","000000000000001110","000000000000011000","111111111111101001","111111111111111011","111111111111111011","000000000000100110","000000000000000100","000000000000101011","111111111111111110","000000000000011101","111111111111101011","000000000000000100","000000000000001010","111111111111110100","000000000000000000","000000000000000010","000000000000011010","000000000000010100","111111111111000010","111111111111111010","000000000000010101","000000000000000001","111111111111110011","000000000000100010","111111111111101001","111111111111101100","000000000000000001","111111111111101101","000000000000011011","111111111111101100","111111111111110111","111111111111101010"),
("111111111111010110","000000000000001110","111111111111001011","000000000000010011","111111111111001010","000000000000000001","000000000000010100","000000000000100010","000000000000010111","000000000000000001","000000000000000001","000000000000010010","111111111111100110","111111111111001101","000000000000000111","000000000000000110","000000000000000111","000000000000001111","111111111111101010","000000000000100110","111111111111100011","111111111111111100","111111111111101111","111111111111110001","111111111111110111","000000000000000011","000000000000000111","000000000000001111","000000000000010010","111111111111111110","000000000000011000","000000000000011011","000000000000100011","000000000000000110","000000000000000111","111111111111111101","111111111111110110","000000000000110001","000000000000010000","000000000000011011","000000000000000100","111111111111101111","000000000000001001","111111111111101101","000000000000001010","111111111111111010","000000000000001110","000000000000100000","000000000000001000","111111111111110001","000000000000000111","000000000000100111","111111111111101110","111111111111111000","000000000000100011","111111111111101100","000000000000010010","000000000000010110","000000000000000011","000000000000001100","000000000000010100","000000000000100101","000000000000010111","111111111111100101","111111111111001111","111111111111111101","111111111111100100","000000000000010001","111111111110110010","111111111111110010","000000000000010001","000000000000010001","000000000000000001","000000000000011111","111111111111111111","000000000000001111","111111111111110101","000000000000110111","111111111111101001","000000000000000101","111111111111101000","000000000000001011","000000000000001111","000000000000001100","000000000000110010","111111111111101000","000000000000000000","000000000000000100","111111111111110001","000000000000000111","000000000000001011","000000000000001100","000000000000100000","111111111111101110","111111111111111111","000000000000000000","000000000000011101","000000000000000111","111111111111100011","000000000000010000","000000000000000101","000000000000001110","000000000000001111","000000000000011010","111111111111101010","000000000000100111","111111111111011110","000000000000001101","000000000000001110","111111111111011000","111111111111110001","000000000000000101","000000000000001000","111111111111111111","111111111111011001","000000000000000001","111111111111111101","000000000000000010","111111111111111100","000000000000100000","000000000000001000","111111111111100110","111111111111110001","111111111111010111","111111111111110010","111111111111010010","111111111111111110","111111111111101111"),
("111111111111110011","000000000000011000","111111111110111010","000000000000001001","111111111110100001","000000000000000110","000000000000000000","000000000000011011","000000000000010111","000000000000010110","111111111111111101","111111111111110010","111111111111101111","111111111111000100","000000000000011010","111111111111110110","000000000000010000","000000000000101001","111111111111111011","000000000000010011","111111111111101111","111111111111011111","111111111111110000","111111111111110000","111111111111101110","000000000000100111","000000000000001111","000000000000011110","000000000000001101","111111111111101100","000000000000100110","111111111111111111","000000000000010111","111111111111100101","111111111111110101","000000000000000010","111111111111100000","000000000000010000","000000000000100000","000000000000001101","000000000000000000","111111111111111010","000000000000000000","000000000000000010","000000000000100111","000000000000001101","000000000000000101","000000000000000010","111111111111110101","111111111111110010","000000000000100101","000000000000100000","000000000000010011","111111111111111111","000000000000011011","111111111111111110","000000000000001011","000000000000001110","111111111111101110","000000000000001010","000000000000000111","000000000000010111","000000000000100110","111111111111101110","111111111111100010","111111111111111110","111111111111000110","000000000000000001","111111111110100110","000000000000000111","000000000000011111","000000000000101110","111111111111111010","000000000000101001","000000000000001101","111111111111111100","111111111111111011","000000000000100000","111111111111101101","111111111111111001","111111111111111000","000000000000000110","111111111111111111","111111111111100001","000000000000101101","111111111111110111","111111111111111010","000000000000001011","111111111111011110","000000000000001010","000000000000011101","000000000000010011","000000000000011101","111111111111101001","000000000000001000","111111111111110110","000000000000011010","000000000000001100","111111111111011110","000000000000001011","111111111111111011","000000000000010001","000000000000000000","000000000000100101","111111111111111111","000000000000001100","000000000000000111","000000000000001110","000000000000000111","111111111111011010","000000000000011000","111111111111110110","000000000000010011","000000000000000010","111111111111001011","000000000000000101","000000000000000001","111111111111111100","111111111111111000","000000000000011101","111111111111100101","000000000000010001","000000000000001101","111111111111001110","000000000000000110","111111111111111000","111111111111110110","000000000000001010"),
("111111111111110001","000000000000010000","111111111110111110","000000000000011111","111111111110100001","000000000000000000","111111111111111000","111111111111111001","000000000000011010","000000000000010011","111111111111110100","111111111111010010","111111111111101100","111111111111010010","111111111111111111","111111111111101011","000000000000010101","000000000000011111","111111111111111110","000000000000011001","111111111111110101","000000000000000110","000000000000010000","111111111111100000","111111111111100011","000000000000000111","111111111111111101","000000000000010010","000000000000011110","111111111111111000","000000000000000000","000000000000000100","111111111111101101","111111111111110101","111111111111111000","000000000000000111","111111111111011011","000000000000001100","000000000000010001","000000000000000001","000000000000001110","111111111111110111","000000000000001011","111111111111101110","000000000000000100","000000000000010011","111111111111111111","000000000000000011","000000000000000000","000000000000000110","000000000000010001","000000000000001110","000000000000010111","111111111111110100","000000000000010101","111111111111101011","000000000000010001","000000000000000110","111111111111110100","111111111111110000","000000000000000000","111111111111111000","000000000000010111","000000000000010011","000000000000001101","000000000000000001","111111111111100000","111111111111110100","111111111110101111","000000000000001111","000000000000010010","000000000000001110","111111111111010110","000000000000010001","000000000000000000","111111111111100111","000000000000000000","000000000000010111","111111111111111000","111111111111110111","111111111111011111","000000000000000000","111111111111111000","111111111111000010","000000000000101100","111111111111111100","111111111111101100","111111111111111011","111111111111100011","000000000000011110","000000000000100110","111111111111101111","000000000000010000","000000000000100100","111111111111100101","111111111111111000","000000000000101001","111111111111100110","111111111111110000","000000000000000001","000000000000001110","000000000000000011","000000000000010011","000000000000101010","111111111111110111","000000000000001111","000000000000000000","111111111111111001","000000000000000000","111111111111110011","111111111111110000","111111111111110101","000000000000010011","111111111111110100","111111111111001000","000000000000010011","111111111111101110","000000000000000101","111111111111101101","111111111111111011","111111111111101010","000000000000011100","000000000000010000","111111111111101001","000000000000001101","111111111111111010","111111111111110011","111111111111110010"),
("111111111111100001","111111111111110100","111111111110111100","000000000000100010","111111111110010001","000000000000001001","111111111111100011","111111111111100100","000000000000010001","000000000000001111","111111111111111110","111111111111110110","111111111111110110","111111111111010001","000000000000001101","111111111111111001","111111111111110100","000000000000001101","111111111111101000","111111111111111101","000000000000000000","111111111111100101","000000000000010101","111111111111100101","111111111111100001","000000000000011010","111111111111100001","000000000000000101","111111111111111010","111111111111010011","111111111111111101","000000000000001100","000000000000000011","111111111111110111","000000000000000111","000000000000010001","111111111111100000","000000000000011101","000000000000000001","111111111111101010","000000000000010000","000000000000001101","111111111111100010","000000000000000100","000000000000001111","000000000000011010","111111111111110000","000000000000000011","111111111111110111","000000000000000001","000000000000000100","000000000000001101","000000000000001010","111111111111100110","000000000000010111","111111111111011010","000000000000100001","000000000000000000","000000000000001010","000000000000000000","000000000000010010","111111111111111101","000000000000000111","000000000000000101","111111111111100101","111111111111101110","111111111111100011","000000000000010011","111111111110110010","000000000000011001","000000000000011100","000000000000010100","111111111111100000","000000000000001101","111111111111111100","111111111111110101","111111111111111111","000000000000101001","111111111111111110","111111111111111101","111111111111100010","000000000000000010","000000000000010100","111111111111001100","000000000000010001","111111111111110011","111111111111110111","000000000000000000","111111111111110000","111111111111111001","000000000000100110","000000000000010100","000000000000011110","000000000000010110","111111111111101011","000000000000010011","000000000000000010","111111111111011110","000000000000000011","111111111111100101","000000000000010100","000000000000000010","111111111111101111","000000000000010110","000000000000001101","000000000000000001","111111111111111110","111111111111110110","111111111111001010","111111111111110100","111111111111110100","000000000000001011","000000000000000001","111111111111110100","111111111111010110","000000000000010000","000000000000010010","111111111111111111","111111111111101011","111111111111110111","111111111111110110","000000000000000000","000000000000011011","111111111111011001","111111111111100101","000000000000010011","111111111111111001","000000000000001000"),
("111111111111011111","000000000000000010","111111111111001011","000000000000011111","111111111111011001","000000000000001010","111111111111111101","111111111111101111","000000000000011100","000000000000001011","111111111111100100","111111111111101111","111111111111011000","111111111111011111","111111111111101000","111111111111101101","000000000000000000","000000000000100001","000000000000000110","000000000000011011","111111111111101110","111111111111011011","000000000000010010","111111111111101000","111111111111101100","000000000000000110","111111111111111110","111111111111111000","111111111111110001","000000000000000000","000000000000001101","000000000000000011","000000000000001101","000000000000101110","111111111111111100","000000000000100100","000000000000000011","000000000000100001","111111111111101010","000000000000010000","000000000000100001","000000000000000100","111111111111011011","000000000000000000","000000000000000000","000000000000011000","111111111111100000","000000000000011110","000000000000000100","111111111111101000","000000000000001001","000000000000000010","000000000000000011","111111111111100001","000000000000010010","111111111111110011","000000000000011010","000000000000001111","111111111111110011","111111111111101110","000000000000000110","000000000000010010","000000000000101101","111111111111110101","111111111111011111","111111111111101111","000000000000000000","000000000000010011","111111111111011001","000000000000100010","000000000000010100","000000000000011000","111111111111100001","111111111111101101","000000000000100011","111111111111100101","111111111111111001","000000000000001001","111111111111010010","111111111111111110","111111111111111101","000000000000000101","111111111111101100","111111111111010111","000000000000101001","000000000000000111","000000000000010001","000000000000000001","000000000000000000","111111111111110100","000000000000010011","000000000000001111","000000000000011101","000000000000100100","111111111111111100","000000000000010001","000000000000011100","111111111111111011","111111111111111111","000000000000000000","000000000000001011","000000000000001001","111111111111110101","000000000000010100","111111111111101011","000000000000011110","111111111111111100","111111111111010101","111111111111001111","111111111111101101","111111111111110100","000000000000011011","000000000000010100","000000000000001001","111111111111100010","000000000000110010","111111111111111100","000000000000000010","111111111111111111","000000000000010000","111111111111111100","000000000000000100","111111111111111110","111111111111101110","111111111111010001","000000000000000100","111111111111100011","000000000000010010"),
("111111111111100001","000000000000010101","111111111111110101","000000000000110110","111111111111110101","000000000000001101","000000000000010010","111111111111111110","000000000000011000","000000000000100010","111111111111111110","111111111111110010","111111111111100011","111111111111110000","111111111111011101","111111111111111011","000000000000001001","000000000000010000","111111111111111001","000000000000000111","111111111111011110","111111111111101010","000000000000001101","111111111111111000","111111111111101101","000000000000000100","111111111111111010","111111111111111001","000000000000000111","111111111111110000","111111111111111001","111111111111110100","000000000000000100","000000000000010011","000000000000010010","000000000000101100","111111111111111100","000000000000101110","111111111111100110","111111111111111101","000000000000000001","000000000000011100","111111111111010111","111111111111101100","000000000000001111","000000000000011110","111111111111011111","000000000000001011","000000000000001001","000000000000000001","111111111111111101","000000000000100010","111111111111110111","111111111111100110","000000000000001000","111111111111010101","000000000000010100","111111111111110001","111111111111110110","111111111111110000","111111111111111110","000000000000010111","000000000000010011","000000000000001000","111111111111100100","111111111111111001","111111111111100100","000000000000001110","111111111111001100","111111111111110001","000000000000010100","000000000000011101","111111111111001101","111111111111011010","000000000000010001","111111111111100010","111111111111111001","000000000000100000","111111111111101000","111111111111110100","111111111111100011","000000000000000101","111111111111111100","111111111111011100","000000000000110010","111111111111011100","000000000000001000","111111111111110111","000000000000001111","111111111111110110","000000000000000111","000000000000011001","000000000000010011","000000000000000111","111111111111101001","000000000000011101","000000000000001001","111111111111101111","111111111111111100","000000000000010000","000000000000001001","000000000000010110","000000000000011001","000000000000110011","111111111111111001","000000000000010100","111111111111110010","111111111111100100","000000000000000000","111111111111110011","000000000000000010","000000000000001110","000000000000011110","000000000000000000","111111111111111010","000000000000100101","000000000000000101","111111111111111001","000000000000000000","111111111111111001","111111111111101101","111111111111100110","111111111111100010","111111111111100110","111111111111110011","000000000000100111","111111111111101101","000000000000000010"),
("000000000000000010","000000000000001000","111111111111111111","000000000000001111","000000000000010110","000000000000010001","000000000000010100","111111111111100100","000000000000000101","000000000000011111","000000000000000100","111111111111100101","111111111111100010","111111111111011010","111111111111001000","000000000000001111","000000000000000011","000000000000101110","000000000000001111","000000000000100001","111111111111011110","111111111111101001","000000000000001000","111111111111110100","111111111111111101","000000000000100000","111111111111010001","111111111111101111","111111111111110100","111111111111100010","000000000000000011","000000000000000000","000000000000101000","000000000000001001","000000000000011100","000000000000011110","000000000000001110","000000000000011010","000000000000000010","000000000000010000","000000000000001101","000000000000011010","111111111110110101","111111111111101011","000000000000001000","000000000000000101","111111111111011110","000000000000010111","111111111111111000","000000000000001001","111111111111111001","000000000000101010","111111111111110000","111111111111111010","111111111111110010","111111111111011100","000000000000000101","000000000000010011","000000000000001111","111111111111110000","000000000000010101","000000000000010001","000000000000100001","000000000000001100","111111111111111111","000000000000011010","111111111111110000","000000000000100010","111111111111110010","111111111111111011","000000000000001001","000000000000000001","111111111111110010","111111111111000110","000000000000001111","000000000000000101","000000000000010010","000000000000000011","111111111111100011","111111111111110011","111111111111101000","000000000000010001","000000000000000001","111111111111010100","000000000000001101","111111111111111000","111111111111111101","000000000000001100","000000000000001010","000000000000000001","000000000000000101","000000000000011011","111111111111101000","000000000000100000","000000000000000011","000000000000000010","111111111111100011","000000000000011001","000000000000000001","111111111111110110","111111111111111110","000000000000000100","000000000000010110","000000000000101111","111111111111101010","000000000000001101","000000000000001100","000000000000001011","111111111111011010","000000000000010001","000000000000000100","000000000000000000","000000000000001110","111111111111111110","000000000000010111","000000000000110010","000000000000000111","111111111111110110","111111111111111001","111111111111101010","000000000000010110","111111111111100110","111111111111100111","111111111111100111","111111111111101011","000000000000100110","000000000000010011","111111111111110110"),
("111111111111111000","000000000000010110","111111111111101110","000000000000011000","000000000000000111","111111111111111001","000000000000001001","111111111111010100","000000000000010001","000000000000010111","111111111111110001","111111111111101001","111111111111100010","111111111111101111","111111111111010101","000000000000001100","000000000000001000","000000000000011010","111111111111111001","000000000000100100","111111111111110100","111111111111100111","000000000000010001","111111111111100111","111111111111101011","000000000000001100","111111111111110110","111111111111011011","000000000000000000","000000000000000111","000000000000010001","111111111111111001","000000000000010001","000000000000011111","000000000000001101","111111111111111011","111111111111111000","000000000000000101","000000000000000000","000000000000011010","000000000000001010","111111111111111010","111111111110111011","111111111111101111","000000000000010011","111111111111111111","111111111111011000","000000000000011011","111111111111111010","111111111111110110","111111111111100110","000000000000100001","000000000000001101","000000000000010011","111111111111111110","111111111111010101","111111111111111000","111111111111110010","000000000000000011","111111111111101110","000000000000000001","000000000000110000","111111111111111010","111111111111101011","000000000000000000","000000000000001001","111111111111110111","000000000000010101","111111111111110001","000000000000000110","111111111111111111","000000000000010110","000000000000001011","111111111111000001","111111111111111111","111111111111110101","000000000000000011","000000000000100000","111111111111010111","000000000000000100","111111111111110101","000000000000011011","111111111111111110","111111111111110100","000000000000101010","111111111111111001","000000000000010010","000000000000011100","111111111111111110","111111111111110010","000000000000001011","000000000000000111","111111111111101101","111111111111111111","111111111111010110","000000000000100001","111111111111101010","000000000000001110","111111111111111110","000000000000000101","000000000000100010","111111111111110110","000000000000101001","000000000000011011","111111111111110101","000000000000010110","000000000000000000","111111111111110011","111111111111111011","000000000000000100","111111111111111101","000000000000010011","000000000000001111","111111111111111101","000000000000101010","000000000000000111","000000000000010111","000000000000010001","111111111111110010","000000000000001001","000000000000001101","000000000000000011","111111111111011011","111111111111110111","111111111111110111","000000000000011000","000000000000000000","000000000000001110"),
("111111111111100100","000000000000001011","111111111111111111","000000000000000110","000000000001000001","000000000000000000","111111111111100010","111111111111101111","111111111111111010","111111111111110011","000000000000000100","111111111111111101","000000000000000101","111111111111101000","111111111111101010","000000000000100100","000000000000001101","000000000000000001","000000000000010001","000000000000010011","111111111111110000","000000000000010001","000000000000011011","000000000000000000","111111111111110110","000000000000000010","000000000000001011","111111111111011010","111111111111111011","111111111111110101","111111111111110111","111111111111101010","111111111111101110","000000000000010010","111111111111111011","000000000000100000","111111111111110010","000000000000001010","111111111111101111","000000000000010000","111111111111110111","000000000000011100","111111111111100101","111111111111110101","000000000000011001","111111111111110101","111111111111110100","000000000000001011","000000000000011011","000000000000000101","111111111111111101","000000000000001010","111111111111101110","000000000000001000","111111111111111011","000000000000000100","111111111111101101","111111111111101100","111111111111110100","111111111111110010","000000000000001011","000000000000001101","000000000000001010","000000000000011001","000000000000001100","000000000000010101","111111111111110110","000000000000001000","111111111111101001","000000000000010111","000000000000000110","000000000000000000","111111111111100100","111111111110101010","000000000000100011","000000000000000000","111111111111111000","111111111111111100","111111111111100001","000000000000000101","000000000000001101","000000000000010000","111111111111110011","000000000000010011","000000000000000100","000000000000000000","111111111111111101","000000000000011011","000000000000001000","111111111111100100","000000000000000000","111111111111110111","111111111111110101","111111111111100111","111111111111000111","000000000000000011","111111111111000000","000000000000000010","000000000000010101","000000000000001111","000000000000010101","000000000000100100","000000000000100100","000000000000010111","111111111111111001","111111111111111111","111111111111111011","000000000000001011","111111111111111101","111111111111111100","111111111111111100","000000000000000000","000000000000000010","111111111111110010","000000000000000111","111111111111111010","000000000000011001","111111111111101011","111111111111011100","000000000000000111","111111111111111101","111111111111101100","111111111111100100","000000000000010011","000000000000000110","000000000000100010","000000000000001010","000000000000001001"),
("000000000000000100","000000000000101010","111111111111111001","000000000000000101","000000000000100110","000000000000000110","111111111111111111","000000000000000000","111111111111111001","000000000000001101","000000000000010000","111111111111110011","111111111111101101","111111111111100100","111111111111011011","111111111111111010","000000000000001101","000000000000000000","000000000000000011","111111111111111100","111111111111001011","000000000000001001","000000000000100101","111111111111110101","111111111111100110","111111111111111110","000000000000011110","111111111111111000","000000000000001100","000000000000000000","111111111111110100","111111111111111010","111111111111111100","000000000000011100","000000000000001011","000000000000001101","111111111111111000","111111111111111110","111111111111101000","111111111111111111","111111111111110111","111111111111111111","111111111111101011","111111111111111111","000000000000011101","111111111111101000","111111111111111111","111111111111111100","111111111111111111","111111111111110011","000000000000000000","000000000000001100","000000000000000000","000000000000001101","000000000000000000","000000000000000010","111111111111101011","111111111111110100","000000000000010111","000000000000000100","000000000000000011","000000000000011001","111111111111110101","000000000000000111","111111111111010001","111111111111111000","111111111111111101","000000000000001111","111111111111111101","000000000000010111","111111111111111000","111111111111101100","111111111111101110","111111111111000010","000000000000000000","111111111111101001","000000000000000010","111111111111101000","111111111111101011","111111111111111100","111111111111111111","000000000000000000","000000000000000111","111111111111110111","000000000000001010","111111111111110100","000000000000010011","000000000000010111","000000000000000001","111111111111100001","111111111111101010","000000000000000111","111111111111100111","111111111111110101","111111111111111011","111111111111110011","111111111111000101","000000000000000111","000000000000000011","000000000000010001","000000000000011001","000000000000001110","000000000000010110","000000000000010110","111111111111110100","000000000000000000","111111111111110011","111111111111011101","111111111111111110","000000000000001010","000000000000000101","000000000000010001","000000000000001111","111111111111110101","000000000000010011","111111111111111111","000000000000010000","111111111111100101","111111111111110010","111111111111111100","000000000000010110","111111111111110000","111111111111001011","000000000000001000","111111111111111111","000000000000100000","000000000000011000","111111111111111101"),
("111111111111110100","000000000000101101","111111111111111111","111111111111011100","000000000000100100","000000000000001111","111111111111111000","000000000000011111","111111111111001100","111111111111100110","111111111111101100","111111111111110001","111111111111101010","111111111111111101","111111111111101011","111111111111111101","000000000000001011","111111111111110100","000000000000100110","000000000000000111","111111111111100110","111111111111111111","000000000000000011","111111111111110011","000000000000000100","111111111111111110","000000000000000011","111111111111011110","111111111111110000","000000000000001010","111111111111101111","111111111111101010","111111111111110011","000000000000010000","000000000000000111","111111111111111111","111111111111111010","000000000000001010","000000000000010001","000000000000000001","000000000000000000","000000000000001000","111111111111110100","111111111111101110","000000000000010110","000000000000001001","000000000000001101","000000000000100101","000000000000110011","000000000000010100","111111111111011000","111111111111110001","111111111111100010","111111111111111000","111111111111101100","111111111111111001","000000000000001101","111111111111110101","000000000000000000","000000000000001000","111111111111110111","111111111111111011","111111111111110010","000000000000000010","111111111110111010","000000000000100010","000000000000010111","000000000000000111","000000000000000111","000000000000010001","111111111111101011","111111111111111110","111111111111110011","111111111111101111","000000000000100001","111111111111011011","111111111111111100","111111111111101101","000000000000000001","111111111111110011","000000000000011100","111111111111111011","111111111111101010","000000000000010100","111111111111101000","111111111111110001","000000000000100100","000000000000001000","000000000000010011","111111111111110001","000000000000001101","000000000000000000","111111111111111011","111111111111011111","111111111111111101","000000000000000000","111111111111100001","111111111111111111","000000000000100001","000000000000011000","111111111111111111","000000000000010011","111111111111110111","000000000000000101","111111111111110110","111111111111101111","111111111111110010","111111111111011000","111111111111110100","000000000000000100","111111111111101010","000000000000000011","000000000000001110","000000000000010101","000000000000011100","111111111111010111","111111111111111111","000000000000000110","111111111111011000","111111111111110111","000000000000010001","000000000000001100","111111111111001100","111111111111111001","111111111111101111","000000000000100000","111111111111101111","000000000000001011"),
("111111111111111000","000000000000100100","000000000000010101","111111111111101101","000000000000100011","000000000000001010","111111111111100111","000000000000011110","111111111111111100","111111111111111001","111111111111111111","000000000000000010","000000000000000111","111111111111100001","111111111111110011","111111111111110010","000000000000010011","111111111111100101","000000000000100110","111111111111110000","111111111111101100","000000000000010101","000000000000100001","000000000000001011","000000000000001100","111111111111101010","000000000000000111","111111111111111000","000000000000010001","111111111111101100","000000000000001001","111111111111111001","000000000000010010","000000000000010010","000000000000001000","111111111111111000","111111111111111100","111111111111110101","000000000000010010","111111111111111110","000000000000101001","000000000000001001","111111111111011100","111111111111101111","000000000000000010","000000000000010101","111111111111101011","111111111111110100","000000000000010101","000000000000010110","111111111111110110","111111111111111110","111111111111110110","000000000000010011","000000000000000000","000000000000000111","000000000000010100","111111111111111111","000000000000001111","111111111111111001","111111111111111000","111111111111110011","111111111111100001","000000000000001010","111111111110100000","000000000000011000","000000000000001101","111111111111111011","000000000000011111","000000000000010110","111111111111100101","111111111111100111","111111111111101111","111111111111100010","000000000000000111","111111111111011100","000000000000000101","111111111111111011","000000000000010011","000000000000001000","000000000000100101","000000000000000110","000000000000001111","000000000000001111","000000000000001100","000000000000010011","000000000000000001","111111111111110100","000000000000000101","111111111111110111","111111111111111011","000000000000001101","111111111111110101","111111111111110010","000000000000010011","000000000000010100","111111111111010101","000000000000000100","111111111111111011","000000000000100000","000000000000001010","111111111111111110","000000000000001001","111111111111111101","111111111111100001","000000000000001010","000000000000000010","111111111111001110","111111111111111010","000000000000100001","000000000000000010","000000000000001010","000000000000000110","000000000000010011","000000000000011110","111111111111100000","000000000000000110","000000000000011001","111111111111110000","000000000000001011","000000000000000010","111111111111101111","111111111111000011","111111111111110111","000000000000001011","000000000000000100","000000000000001000","111111111111100100"),
("000000000000011110","111111111111111100","000000000000000000","111111111111010001","000000000000001100","000000000000001001","000000000000000000","000000000000011001","111111111111010011","111111111111011100","111111111111111111","000000000000011000","111111111111111011","111111111111111100","111111111111101001","111111111111010001","111111111111101001","111111111111110101","000000000000011100","111111111111001100","111111111111101110","000000000000010010","000000000000000001","111111111111110100","000000000000000110","000000000000001100","000000000000000000","111111111111101110","111111111111110111","111111111111111100","000000000000000000","111111111111011111","000000000000000010","000000000000011011","000000000000101100","111111111111110011","000000000000011011","111111111111111111","000000000000011110","000000000000000000","000000000000011101","000000000000010111","111111111111110111","111111111111101111","000000000000001100","000000000000000110","111111111111101100","000000000000110111","000000000000100000","000000000000000101","111111111111110000","111111111111110100","000000000000000000","000000000000000000","111111111111100111","000000000000000000","000000000000001010","111111111111001101","000000000000000110","111111111111110011","111111111111101101","111111111111100101","111111111111001001","000000000000000111","111111111110111111","000000000000010111","000000000000011000","000000000000000000","000000000000011011","111111111111111101","111111111111100010","111111111111011011","000000000000100001","111111111111101111","000000000000000101","111111111111100001","000000000000010111","111111111111110110","000000000000001110","111111111111111101","000000000000111011","000000000000000011","111111111111111101","111111111111111101","111111111111011111","000000000000001110","000000000000000110","000000000000001111","000000000000010111","111111111111011101","000000000000000110","000000000000000111","111111111111100000","111111111111100100","000000000000011000","000000000000000010","111111111111111100","111111111111111001","000000000000001000","000000000000001101","000000000000011000","000000000000011100","000000000000010010","111111111111110010","111111111111110010","111111111111110111","000000000000010111","111111111111101000","000000000000000001","000000000000011010","111111111111100011","111111111111111110","000000000000010010","111111111111110001","000000000000101110","111111111111101000","111111111111101100","000000000000010100","000000000000001000","111111111111100100","000000000000010010","000000000000101101","111111111111010011","000000000000000110","000000000000001001","111111111111011100","000000000000000101","111111111111100010"),
("111111111111110101","111111111111001001","000000000000010110","111111111111100000","111111111111001011","000000000000000101","111111111111110010","000000000000001010","111111111111111001","111111111111000001","111111111111011101","000000000000100001","000000000000011100","111111111111101111","000000000000000001","111111111111011001","111111111111110111","111111111111111001","000000000000001110","000000000000000011","111111111111010100","111111111111110100","111111111111010101","111111111111101100","000000000000010001","000000000000000110","111111111111110100","111111111111101010","000000000000010000","111111111111110001","000000000000010010","111111111111101100","000000000000010110","111111111111101011","000000000000011101","000000000000000110","000000000000100000","111111111111111101","000000000000010110","000000000000010101","000000000000100110","000000000000101101","111111111111111101","111111111111010101","000000000001000010","111111111111111101","111111111111101011","000000000000101010","000000000000101000","000000000000000111","111111111111110101","000000000000010010","000000000000001011","000000000000001101","000000000000000100","000000000000000000","000000000000100010","111111111111101011","000000000000000000","111111111111111001","000000000000000100","111111111111011101","111111111111001011","111111111111111110","111111111111100010","000000000000110101","000000000000011001","111111111111110101","000000000000100110","000000000000011001","111111111111111011","111111111111111101","000000000000010010","111111111111110001","111111111111111010","111111111111110011","000000000001000100","111111111111111110","000000000000011011","111111111111111110","000000000000010110","000000000000100110","111111111111100111","111111111111100001","111111111111100101","111111111111111011","000000000000100011","111111111111110111","000000000000001011","000000000000000000","111111111111100011","111111111111101111","111111111111110100","111111111111011100","000000000000011111","000000000000011110","000000000000000011","111111111111101000","111111111111111100","111111111111110111","000000000000000011","000000000000111010","111111111111101001","000000000000000110","000000000000010010","000000000000000110","000000000000011000","111111111111111101","111111111111111100","111111111111110011","000000000000001010","111111111111110001","000000000000010110","000000000000000000","000000000000101100","111111111111011010","111111111111111010","000000000000011110","111111111111101100","111111111111111111","000000000000011000","000000000000000101","111111111111011111","111111111111101101","111111111111110001","111111111111001011","111111111111110100","000000000000010001"),
("000000000000000000","111111111111100111","111111111111110111","000000000000000100","111111111111100000","000000000000000011","111111111111110010","000000000000010111","111111111111111110","111111111111000111","000000000000001010","000000000000111000","000000000000001100","111111111111111101","000000000000000101","111111111111110010","111111111111111010","000000000000000101","000000000000101110","000000000000001111","111111111111110110","000000000000010111","111111111111001110","000000000000001110","000000000000010101","000000000000010011","000000000000000101","111111111111111010","111111111111111101","111111111111101111","000000000000001100","111111111111011111","000000000000101011","000000000000000000","000000000000101010","000000000000000110","000000000000010001","000000000000011001","111111111111110000","111111111111111101","000000000000001101","000000000000010010","000000000000011001","111111111111011111","000000000001000110","111111111111111110","000000000000000100","000000000000101010","000000000000011001","000000000000000100","111111111111100001","000000000000001110","000000000000000101","000000000000100001","000000000000000001","000000000000010110","000000000000101001","111111111111010100","000000000000001101","111111111111111000","000000000000000111","111111111111101100","111111111111100011","111111111111011000","111111111111010001","000000000000100000","000000000000010110","111111111111100111","000000000000100111","000000000000000100","111111111111101100","111111111111110001","111111111111100101","111111111111100111","111111111111100010","111111111111111001","000000000001000000","111111111111110111","000000000000000011","000000000000010011","111111111111110000","000000000000110001","000000000000000101","111111111111101110","111111111111111101","111111111111011011","000000000000001111","000000000000000100","000000000000000101","111111111111111100","000000000000000110","000000000000000010","000000000000001100","111111111111010100","000000000000100001","000000000000011111","000000000000000111","111111111111110110","111111111111101110","000000000000100001","111111111111111010","000000000000110000","111111111111100100","000000000000010100","000000000000100000","000000000000001000","000000000000010011","000000000000000000","111111111111111100","000000000000001100","000000000000000111","000000000000000101","000000000000001000","000000000000001010","000000000000101100","111111111111101001","000000000000000010","000000000000110001","000000000000000011","000000000000000000","000000000000010000","111111111111111100","111111111111110010","111111111111110110","111111111111010001","111111111111111011","000000000000000010","111111111111111010"),
("000000000000100011","111111111111111100","000000000000000000","111111111111111111","111111111111101111","111111111111110001","000000000000000100","000000000000010101","000000000000001010","111111111111100110","111111111111111010","000000000000110101","000000000000010001","111111111111010101","111111111111111110","111111111111111000","111111111111101010","000000000000011111","000000000000011111","000000000000001110","000000000000001000","000000000000000001","111111111111110101","000000000000001001","000000000000101100","111111111111111100","111111111111101000","111111111111111010","111111111111101111","111111111111111010","000000000000010000","111111111111110101","000000000000000010","000000000000000100","111111111111111100","000000000000001111","111111111111110100","111111111111101111","111111111111110111","111111111111100011","000000000000010101","000000000000011101","000000000000101101","111111111111101111","000000000000100110","111111111111110101","000000000000001010","000000000000011010","000000000000010010","000000000000011010","111111111111101100","000000000000000010","000000000000100011","000000000000011001","111111111111111011","000000000000000100","000000000000101110","000000000000011011","000000000000010000","000000000000001010","000000000000100011","111111111111101101","111111111111101101","111111111111111011","111111111111110011","000000000000011100","000000000000000011","000000000000001011","111111111111111001","111111111111101110","000000000000010110","111111111111110101","000000000000011101","111111111111110110","000000000000001011","111111111111110111","000000000000101101","111111111111111101","111111111111100000","000000000000001110","111111111111011110","000000000000101000","111111111111010110","111111111111100011","000000000000001010","111111111111010011","000000000000101100","111111111111110110","111111111111111000","111111111111100010","111111111111110000","000000000000011000","111111111111110000","111111111111001111","000000000000100100","000000000000001111","111111111111110110","000000000000000000","111111111111110111","000000000000010101","000000000000100000","000000000000110100","000000000000100111","000000000000001110","000000000000001110","111111111111111101","000000000000001001","000000000000001100","111111111111101001","000000000000000001","000000000000010110","000000000000001010","000000000000011010","000000000000110000","000000000000000001","000000000000010000","000000000000010010","000000000000101000","111111111111100011","000000000000000100","000000000000110100","111111111111110010","000000000000010100","111111111111111001","111111111111101011","000000000000000000","000000000000001100","000000000000001001"),
("000000000000101000","000000000000001100","111111111111110010","111111111111110010","000000000000000110","000000000000011000","000000000000000111","111111111111110001","111111111111110101","000000000000000000","111111111111110010","000000000000000001","111111111111110000","111111111111011110","000000000000001100","000000000000010110","000000000000000000","111111111111110001","111111111111111001","111111111111100110","000000000000000000","111111111111111101","111111111111111110","111111111111101001","000000000000000000","000000000000010010","111111111111111000","000000000000010000","000000000000010011","000000000000001001","111111111111011110","000000000000000100","000000000000000010","111111111111111101","111111111111111100","111111111111111001","111111111111110110","111111111111111100","111111111111110111","111111111111111011","111111111111101111","111111111111111110","000000000000000101","000000000000001101","000000000000010010","000000000000001000","000000000000101001","111111111111110000","111111111111111000","000000000000011101","111111111111011101","111111111111100111","111111111111111000","000000000000000001","000000000000000011","111111111111110001","111111111111101110","000000000000001000","000000000000000000","111111111111101110","111111111111110000","111111111111111001","111111111111101010","111111111111111101","111111111111111110","000000000000001111","111111111111111101","000000000000100001","000000000000000111","111111111111111111","000000000000010001","111111111111101100","000000000000001110","111111111111110111","000000000000000111","000000000000000111","000000000000000111","111111111111110111","000000000000000111","000000000000010011","000000000000001001","000000000000001001","111111111111111111","111111111111100101","111111111111101000","111111111111101011","111111111111110101","000000000000000001","000000000000001101","000000000000000111","000000000000001010","000000000000010100","111111111111111011","111111111111110110","000000000000000011","000000000000001110","000000000000000010","111111111111110110","000000000000010110","000000000000100011","000000000000000110","000000000000101110","000000000000001000","111111111111100011","111111111111101111","000000000000001010","111111111111111100","000000000000000000","000000000000000000","000000000000010011","000000000000001010","111111111111111110","000000000000010101","000000000000000011","111111111111010011","000000000000100110","000000000000010000","000000000000000010","000000000000000000","111111111111111010","000000000000001111","111111111111100111","111111111111110111","111111111111110111","000000000000001100","000000000000010010","000000000000011010","000000000000001101"),
("111111111111110001","000000000000001101","111111111111101111","111111111111101111","111111111111101100","000000000000000000","000000000000001111","111111111111111001","111111111111111101","000000000000001101","111111111111101100","111111111111101101","111111111111110110","000000000000000100","111111111111111001","111111111111110100","000000000000000000","111111111111111000","111111111111110101","000000000000000111","111111111111101100","000000000000010010","000000000000001001","000000000000010000","111111111111110101","000000000000000101","000000000000001011","111111111111111011","000000000000001110","111111111111101111","111111111111110010","111111111111111111","111111111111111001","000000000000001011","111111111111110001","000000000000010011","000000000000010100","000000000000001011","111111111111111101","111111111111111101","111111111111101111","000000000000000001","111111111111101101","000000000000001011","000000000000001001","111111111111111000","000000000000001000","111111111111111011","000000000000000000","000000000000001011","111111111111101101","000000000000000001","111111111111111001","111111111111101100","000000000000000000","111111111111111101","000000000000000101","000000000000000000","000000000000001000","111111111111111000","111111111111110110","000000000000000110","111111111111110000","111111111111110011","000000000000000010","111111111111110000","000000000000000110","111111111111111000","111111111111101101","111111111111110000","000000000000010000","111111111111110100","000000000000001010","111111111111110111","111111111111111001","111111111111110110","111111111111111010","111111111111110100","000000000000010010","000000000000010000","000000000000001101","000000000000000001","111111111111110011","000000000000000000","111111111111110001","111111111111110111","000000000000001101","000000000000000000","000000000000001010","000000000000010001","000000000000001010","000000000000000000","111111111111110110","000000000000010001","111111111111110011","000000000000000001","111111111111110001","000000000000000000","000000000000001100","000000000000000000","000000000000001110","111111111111101101","000000000000010001","000000000000001100","111111111111111110","111111111111110000","111111111111101110","111111111111111001","000000000000000100","000000000000001101","000000000000001111","111111111111111011","000000000000000000","000000000000000010","111111111111101101","000000000000000000","111111111111111011","000000000000000000","111111111111111111","000000000000001010","000000000000001011","000000000000001111","000000000000001101","111111111111101111","111111111111111100","000000000000000011","111111111111110010","000000000000000100"),
("000000000000010000","111111111111111100","000000000000001100","111111111111111111","111111111111101111","000000000000001010","111111111111101100","111111111111110001","111111111111110011","111111111111111011","000000000000010010","111111111111111111","000000000000000100","111111111111111000","000000000000000011","000000000000000101","000000000000000101","000000000000001000","111111111111101111","111111111111101111","000000000000010011","111111111111110000","000000000000000000","000000000000001000","000000000000000000","000000000000000110","111111111111110110","111111111111111110","111111111111111000","111111111111111100","000000000000000101","000000000000010000","111111111111110000","111111111111101101","000000000000000001","000000000000000100","000000000000001101","111111111111110100","000000000000001000","111111111111111100","111111111111101110","111111111111110001","000000000000010010","111111111111110011","000000000000010001","111111111111111110","000000000000001110","111111111111101111","000000000000001000","111111111111110100","111111111111110101","111111111111110011","000000000000001011","000000000000010001","111111111111111101","000000000000010100","000000000000000011","000000000000001001","111111111111111110","000000000000001110","111111111111111010","000000000000010010","111111111111110011","111111111111110010","000000000000001011","111111111111101110","111111111111111000","000000000000000010","000000000000000000","111111111111101110","111111111111110010","111111111111101111","000000000000000110","111111111111111011","111111111111111011","111111111111111000","000000000000000000","000000000000010100","111111111111110111","000000000000000000","000000000000000100","000000000000001010","000000000000001000","000000000000001000","111111111111110001","000000000000010001","000000000000000110","000000000000000000","111111111111110110","111111111111111111","111111111111110011","111111111111111010","000000000000000001","111111111111101101","111111111111110010","000000000000000000","000000000000001100","111111111111110010","111111111111111001","111111111111101100","000000000000000101","111111111111110110","000000000000000000","000000000000000101","111111111111111110","000000000000010001","000000000000001101","000000000000010000","111111111111110001","000000000000010011","111111111111110110","111111111111111011","111111111111111001","111111111111111000","111111111111110001","111111111111111011","000000000000001101","000000000000000000","111111111111101101","000000000000010010","111111111111111001","000000000000000111","000000000000010100","000000000000000100","111111111111111110","111111111111110011","000000000000000110","111111111111110101"),
("111111111111111000","111111111111101110","111111111111101011","000000000000101110","000000000000000010","000000000000010011","111111111111111001","000000000000000010","000000000000101001","000000000000000010","000000000000010001","000000000000000101","000000000000100100","000000000000100101","000000000000000000","000000000000000110","111111111111101111","000000000000000110","000000000000001110","000000000000000000","000000000000000101","111111111111100010","000000000000001011","000000000000010110","000000000000000001","000000000000001000","000000000000001101","000000000000010001","000000000000010101","111111111111111101","000000000000000000","000000000000001110","111111111111100101","111111111111110100","111111111111101111","000000000000101101","111111111111110010","111111111111111101","000000000000001000","111111111111110100","111111111111101010","000000000000000101","111111111111101000","000000000000001100","111111111111011101","000000000000001010","000000000000001011","000000000000010111","111111111111100010","111111111111110001","111111111111110010","111111111111100111","111111111111111101","111111111111110110","000000000000010110","111111111111101100","111111111111110100","111111111111110111","111111111111010110","111111111111110000","000000000000000110","000000000000010111","000000000000011101","000000000000011001","000000000000110100","111111111111111000","000000000000000110","111111111111110010","000000000000000001","000000000000001111","000000000000100001","000000000000011000","000000000000000000","111111111111111100","000000000000001111","111111111111110100","111111111111110010","111111111111111001","000000000000000110","111111111111010111","000000000000010101","111111111111110010","111111111111111000","000000000000100010","000000000000100100","000000000000000101","000000000000001001","111111111111111110","111111111111100000","000000000000011111","000000000000000001","111111111111110111","111111111111111111","000000000000100111","111111111111010100","111111111111011011","111111111111110111","000000000000000001","000000000000000100","111111111111100100","111111111111110010","000000000000001010","111111111111111101","000000000000100001","000000000000011001","000000000000011010","000000000000001001","111111111111001100","111111111111110111","111111111111111010","111111111111111111","000000000000000100","111111111111101000","000000000000001011","000000000000001010","000000000000000100","111111111111101100","000000000000010110","000000000000011110","000000000000000111","111111111111101110","000000000000001010","000000000000000011","000000000000001110","111111111111110001","111111111111110010","111111111111111101","000000000000000110"),
("000000000000001010","111111111111111000","111111111111111101","111111111111111100","111111111111100010","000000000000000111","000000000000000111","000000000000000101","000000000000001000","111111111111101100","000000000000001111","111111111111101111","000000000000001111","000000000000000010","111111111111111000","111111111111111011","000000000000000001","000000000000011011","000000000000001011","000000000000000101","111111111111110010","111111111111111011","000000000000000111","000000000000011110","111111111111111111","000000000000001001","000000000000000000","111111111111111010","000000000000010000","000000000000000111","000000000000011111","111111111111110001","000000000000000111","111111111111111000","111111111111100100","111111111111111010","111111111111111000","000000000000001001","111111111111111011","111111111111110110","111111111111110100","111111111111110110","111111111111111011","111111111111110011","111111111111111110","000000000000000100","111111111111101101","000000000000011010","111111111111111000","111111111111011100","111111111111110001","000000000000010011","111111111111111111","111111111111111111","000000000000101001","000000000000011100","111111111111011111","000000000000001100","111111111111110010","000000000000001101","111111111111110101","000000000000001110","111111111111110101","111111111111110111","000000000000000001","111111111111101011","000000000000011110","111111111111100001","111111111111101011","000000000000001101","000000000000001001","000000000000010100","000000000000011010","000000000000010110","111111111111111011","000000000000010000","000000000000001000","000000000000000100","111111111111101111","000000000000010110","000000000000000000","000000000000000001","111111111111110110","000000000000000110","111111111111111101","111111111111001110","111111111111011011","000000000000010110","111111111111111111","000000000000000101","111111111111101000","000000000000001111","111111111111101100","000000000000010001","111111111111101111","000000000000000100","000000000000010001","000000000000001101","000000000000000111","111111111111100100","000000000000010000","111111111111101110","000000000000001000","000000000000011011","000000000000000100","000000000000000100","111111111111101100","111111111111010010","000000000000000000","000000000000001111","111111111111110010","111111111111111001","111111111111111001","111111111111110100","000000000000010101","111111111111110010","000000000000000011","000000000000001000","000000000000000010","111111111111110010","000000000000000011","111111111111111100","111111111111100110","000000000000000000","111111111111111000","111111111111100011","111111111111110110","111111111111111011"),
("111111111111011000","000000000000001010","111111111111100100","111111111111101001","111111111111101111","000000000000101010","000000000000011000","111111111111100111","111111111111111101","000000000000011110","000000000000001100","111111111111100010","000000000000101110","111111111111110011","000000000000101010","000000000000001010","000000000000001110","111111111111101110","000000000000000111","000000000000010010","111111111110111110","111111111111000101","000000000000001000","111111111111101001","111111111111101010","000000000000011110","111111111111010011","111111111111101110","000000000000100001","111111111111100100","000000000000000101","000000000000011101","000000000000001101","111111111111001011","111111111111101000","000000000000001000","000000000000000110","111111111111100001","111111111111111010","111111111111100101","111111111111101100","111111111111010010","000000000000111101","000000000000100000","000000000000000000","000000000000000000","000000000000011111","000000000000000100","111111111111101011","111111111111111000","000000000000001010","000000000000000000","000000000000001100","111111111111101010","000000000000011010","111111111111110001","111111111111011001","000000000000000000","111111111111110111","111111111111110101","000000000000011111","000000000000001111","111111111111110111","000000000000010000","111111111111111010","111111111111011001","000000000000110100","000000000000000111","111111111111101101","000000000000000000","000000000000001011","000000000000000101","000000000000101111","000000000000011111","000000000000011010","000000000000010001","111111111111011101","000000000000010101","111111111111111100","000000000000001110","000000000000000010","111111111111100000","000000000000100111","000000000000000000","000000000000000001","111111111111101000","111111111111010101","000000000000001000","111111111111111010","000000000000101010","111111111111010011","111111111111110001","111111111111101100","111111111111100100","111111111111101111","000000000000001010","000000000000101010","000000000000000101","111111111111010101","000000000000100001","111111111111111110","111111111111101010","000000000000000111","000000000000100010","000000000000001010","000000000000000110","111111111111110100","000000000000011110","111111111111111011","111111111111111101","111111111111101111","000000000000000110","000000000000001000","111111111111101101","111111111111010000","111111111111110101","000000000000101011","111111111111101010","111111111111111010","000000000000001011","111111111111110000","111111111111011001","111111111111101101","000000000000011100","000000000000101000","111111111111100110","000000000000000000","111111111111111100"),
("111111111111101100","000000000000000100","111111111111100000","111111111111110101","000000000000110111","000000000000010100","111111111111110000","111111111111100110","000000000000010101","000000000000010000","111111111111101100","111111111111101001","000000000000101110","111111111111100110","000000000000101010","111111111111100010","111111111111110011","111111111111110111","000000000001000110","000000000000001101","111111111111011111","111111111110111100","000000000000010000","000000000000010100","111111111111011000","111111111111100010","111111111111111010","111111111111100110","000000000000100110","111111111111111010","111111111111101101","000000000000100000","111111111111100100","111111111111011001","111111111111101010","111111111111111010","111111111111111100","000000000000010000","111111111111111010","000000000000000010","000000000000101010","111111111111101000","000000000000001010","000000000000010001","111111111111100100","000000000000000010","000000000000110000","111111111111111100","111111111111111011","000000000000011111","111111111111111001","111111111111111000","000000000000000111","000000000000010010","000000000000100000","000000000000010001","111111111111101001","000000000000010101","000000000000000000","111111111111111011","111111111111111110","000000000000000100","111111111111111010","111111111111111110","111111111111010100","111111111111011100","000000000000010101","111111111111011111","111111111111100100","111111111111101101","000000000000000011","000000000000100110","000000000000110110","000000000000000001","000000000000110010","111111111111111000","111111111111001100","111111111111111001","000000000000001101","000000000000000110","111111111111100100","111111111111001000","000000000000001011","000000000000100010","111111111111111000","111111111111110110","111111111111111100","000000000000010111","111111111111111000","000000000000100110","111111111111011000","111111111111111011","111111111111110010","111111111111101111","111111111111011011","000000000000001011","000000000000101000","111111111111110100","111111111111110000","000000000000001100","000000000000001000","111111111111001110","111111111111101010","000000000000001000","000000000000000100","111111111111011111","000000000000000011","000000000000001110","111111111111111111","000000000000010011","111111111111100110","111111111111110111","111111111111110010","000000000000000111","111111111111011010","111111111111011110","111111111111101111","000000000000010100","111111111111011101","000000000000001011","111111111111111111","111111111111110000","000000000000000000","000000000000000111","000000000000011001","111111111111001011","111111111111101011","000000000000011001"),
("111111111111001011","000000000000001001","111111111111101000","111111111111111011","000000000000110110","000000000000010001","000000000000001010","000000000000000000","000000000000010011","000000000000010100","111111111111111010","000000000000000001","000000000000000111","111111111111000110","000000000000011100","111111111111110010","000000000000000110","111111111111111100","000000000000011010","000000000000001110","111111111110111001","111111111111011011","000000000000000000","000000000000011011","111111111111101010","111111111111101110","000000000000100100","111111111111011011","000000000000100000","111111111111011101","111111111111110100","111111111111111111","111111111111100110","111111111110111111","111111111111101010","000000000000010000","111111111111111110","000000000000001010","111111111111110000","000000000000000010","000000000000101001","111111111111101110","000000000000001011","000000000000000001","111111111111010101","000000000000010001","000000000000001101","000000000000000010","111111111111110110","000000000000001000","000000000000000100","000000000000000010","000000000000000100","111111111111111111","000000000000010111","000000000000001000","111111111111111000","000000000000000100","000000000000001011","111111111111110111","111111111111110011","000000000000001010","000000000000000000","000000000000000100","111111111111011011","111111111111101011","000000000000001011","111111111111101100","111111111111101100","111111111111100100","000000000000010100","000000000000011001","000000000000011101","111111111111111110","000000000000100000","111111111111101111","111111111111101001","111111111111111110","000000000000010011","000000000000000000","111111111111111001","111111111111001101","000000000000100100","000000000000000010","000000000000000010","000000000000000000","111111111111101010","000000000000000001","111111111111100111","000000000000110000","111111111111010101","111111111111110101","111111111111111001","111111111111110110","111111111111101110","111111111111110010","000000000000011001","111111111111101010","111111111111011000","000000000000000100","000000000000010000","111111111111111011","111111111111111000","000000000000000101","111111111111011001","111111111111110000","000000000000001000","000000000000010101","000000000000000011","000000000000000101","111111111111110001","111111111111101010","111111111111011111","000000000000011000","111111111111111000","111111111111101110","000000000000001000","000000000000100011","111111111111111000","000000000000010111","111111111111111000","111111111111011000","000000000000000100","111111111111110110","000000000000101101","111111111111001000","000000000000000001","000000000000000000"),
("111111111111011100","111111111111111100","111111111111101111","111111111111101110","000000000001000000","111111111111110110","111111111111111111","000000000000110001","000000000000010101","000000000000010001","000000000000000011","000000000000000110","000000000000001000","111111111111110000","000000000000011111","000000000000001011","111111111111110101","000000000000001001","000000000000111011","000000000000001101","111111111111100010","111111111111001001","111111111111011111","111111111111111010","111111111111011000","000000000000001000","000000000000100010","111111111111110111","000000000000101001","111111111111011111","111111111111010011","000000000000000001","000000000000000100","111111111110110001","111111111111101000","000000000000010111","111111111111111010","000000000000001011","111111111111111001","000000000000001010","111111111111111010","111111111111011111","000000000000000101","000000000000000000","111111111111101100","000000000000010111","000000000000010000","111111111111100100","000000000000001011","111111111111111100","000000000000100110","111111111111101110","000000000000000111","000000000000001110","111111111111111101","111111111111101011","000000000000000100","000000000000010001","000000000000001010","111111111111110001","111111111111111010","000000000000000001","111111111111111001","000000000000001001","111111111111100100","111111111111100100","000000000000001100","000000000000000011","000000000000000101","111111111111101111","000000000000000100","000000000000101011","000000000000010001","000000000000001100","000000000000000110","111111111111100101","111111111111111101","111111111111101110","000000000000010101","000000000000001010","111111111111110010","111111111111110001","000000000000010100","000000000000010011","000000000000010001","111111111111010111","000000000000000001","111111111111101111","000000000000010000","000000000000011111","111111111111001100","000000000000000101","000000000000000001","111111111111010011","111111111111010101","000000000000000000","000000000000010101","000000000000001101","111111111111100100","000000000000011001","111111111111101101","111111111111110001","000000000000000111","000000000000000010","111111111111110010","111111111111100001","111111111111100000","000000000000011100","000000000000011010","111111111111111100","111111111111101110","111111111111101010","000000000000001010","000000000000001010","000000000000000111","000000000000000011","000000000000010101","000000000000001001","111111111111110001","000000000000000001","000000000000000110","111111111111011000","111111111111111100","111111111111101110","000000000000001101","111111111111101100","111111111111111101","111111111111110101"),
("111111111111000111","000000000000001101","111111111111100001","111111111111111111","000000000000101110","111111111111101100","000000000000000100","111111111111111110","000000000000000010","000000000000001100","111111111111110100","000000000000000100","111111111111100010","111111111111100000","000000000000111100","000000000000000010","000000000000000100","111111111111111110","000000000000010111","000000000000000110","111111111111000100","111111111111110011","111111111111110010","111111111111011000","111111111111011011","111111111111110010","111111111111111011","111111111111111111","000000000000000001","111111111111000101","111111111111011111","111111111111101110","000000000000000000","111111111111101001","111111111111111001","111111111111111111","000000000000100011","111111111111110100","000000000000010000","111111111111110110","111111111111111010","111111111111110110","000000000000011011","000000000000000111","111111111111110100","000000000000000000","000000000000010101","111111111111101001","111111111111111111","111111111111111110","000000000000011101","000000000000000111","000000000000000000","111111111111110101","000000000000010110","111111111111110010","111111111111100010","000000000000011100","000000000000010100","000000000000001110","111111111111111101","000000000000000111","111111111111110001","111111111111111011","111111111111010110","111111111111111111","111111111111110010","000000000000000001","111111111111011101","111111111111011011","111111111111110000","000000000000001111","111111111111110111","000000000000000110","111111111111111001","111111111111100000","000000000000001111","111111111111110100","000000000000011011","000000000000100011","111111111111101010","111111111111100111","111111111111110110","111111111111111010","000000000000000010","111111111111110111","000000000000000010","111111111111111001","000000000000000000","000000000000010010","111111111111010000","111111111111101100","000000000000011001","111111111111101000","111111111111110111","111111111111011011","111111111111111000","000000000000011000","111111111111011010","000000000000001011","111111111111110101","000000000000011001","000000000000000011","111111111111110011","000000000000000110","111111111111100110","111111111111100100","000000000000100011","000000000000000000","000000000000000110","111111111111110110","000000000000001011","111111111111111010","000000000000010100","111111111111100001","111111111111110000","111111111111110111","000000000000000111","111111111111110010","000000000000000100","000000000000001010","111111111111111100","000000000000000010","000000000000010000","000000000000011111","111111111111101011","111111111111111100","111111111111100111"),
("111111111111000101","111111111111110110","111111111111110100","111111111111100001","000000000000101010","111111111111111010","000000000000000011","000000000000000001","000000000000010101","000000000000010011","111111111111111100","000000000000010111","111111111111111010","111111111111100100","000000000000100001","111111111111110100","111111111111111010","000000000000000000","000000000000000000","000000000000011010","111111111111010110","000000000000000111","000000000000001111","111111111111010111","111111111111011100","000000000000000101","000000000000010110","111111111111110111","111111111111110000","111111111111111011","111111111111110110","000000000000000111","111111111111101100","000000000000000101","000000000000010001","111111111111110000","000000000000000001","111111111111110111","111111111111111100","000000000000011001","000000000000001100","000000000000001001","000000000000000101","111111111111100010","000000000000000100","111111111111111000","000000000000001001","000000000000010001","000000000000100000","000000000000001100","000000000000010000","000000000000011000","111111111111111000","111111111111101000","000000000000010001","111111111111101110","111111111111111010","000000000000000110","000000000000011110","000000000000001010","000000000000000100","000000000000001100","000000000000000011","111111111111110100","111111111110110011","000000000000001011","111111111111101111","111111111111101000","111111111111011100","111111111111010111","111111111111110001","000000000000000100","111111111111110001","000000000000010010","111111111111111101","000000000000000100","000000000000001001","111111111111110101","000000000000010110","000000000000011110","111111111111101110","000000000000001010","000000000000010100","000000000000010000","111111111111111111","111111111111101110","000000000000011110","000000000000000101","111111111111111011","000000000000001101","111111111111100100","000000000000000010","000000000000011100","111111111111011001","000000000000001101","111111111111101011","000000000000011001","000000000000101000","111111111110111101","000000000000011110","111111111111100101","000000000000000110","111111111111110000","111111111111111010","111111111111110100","111111111111111010","111111111111111010","111111111111111111","000000000000001111","000000000000000011","000000000000000101","111111111111111011","111111111111111110","111111111111110101","111111111111010111","111111111111110111","000000000000001001","000000000000000000","111111111111110001","000000000000011110","000000000000001001","000000000000000001","000000000000010101","000000000000000000","000000000000010000","000000000000000000","000000000000010010","111111111111100101"),
("111111111111100000","000000000000001010","111111111111001111","111111111111110100","000000000000000110","111111111111100101","111111111111100110","000000000000100111","111111111111101111","111111111111110110","000000000000001010","000000000000010001","111111111111011000","111111111111110100","111111111111111111","000000000000011011","111111111111110001","000000000000010100","111111111111110100","111111111111111110","111111111111001111","000000000000010000","000000000000011000","111111111111011011","111111111111111111","000000000000000000","000000000000001101","000000000000000000","111111111111110010","000000000000000100","111111111111110110","111111111111111110","000000000000001110","111111111111111101","111111111111111101","000000000000000010","000000000000001011","111111111111111000","111111111111111010","000000000000000011","111111111111111010","111111111111111010","111111111111110111","111111111111111001","000000000000000011","000000000000000100","000000000000001010","000000000000001101","000000000000000111","111111111111110101","111111111111110100","111111111111111011","000000000000000010","111111111111100111","000000000000010110","111111111111110101","111111111111101110","000000000000010100","000000000000000101","000000000000001010","111111111111111110","000000000000101010","000000000000001001","111111111111011000","111111111111001001","111111111111110000","111111111111010001","000000000000000011","111111111111100001","111111111111110000","111111111111111101","000000000000000101","000000000000010010","111111111111111000","111111111111111100","111111111111101111","000000000000001101","000000000000001111","000000000000010001","000000000000000000","111111111111111100","000000000000100101","000000000000000011","000000000000000111","000000000000011010","111111111111101010","111111111111111101","000000000000010111","000000000000001101","000000000000010101","000000000000000001","000000000000001101","000000000000111000","111111111111110111","111111111111111100","000000000000000001","000000000000001110","000000000000001000","111111111111100111","000000000000001010","111111111111111110","000000000000010101","000000000000000010","111111111111110111","111111111111111011","111111111111100000","000000000000001010","111111111111110001","000000000000000001","111111111111100010","000000000000001101","000000000000000001","000000000000000011","111111111111110110","111111111111100010","111111111111011110","111111111111110101","111111111111110001","111111111111111101","000000000000101010","000000000000000000","111111111111111101","111111111111111101","000000000000001010","111111111111111000","111111111111101011","000000000000000101","111111111111100111"),
("111111111111101001","000000000000000110","111111111111011001","111111111111110101","111111111110011110","111111111111110111","111111111111110000","000000000000010111","000000000000011110","111111111111111001","111111111111110101","000000000000010110","111111111111010111","111111111111000101","111111111111110110","000000000000010101","000000000000000000","000000000000011100","000000000000000000","111111111111111101","111111111111010011","111111111111101100","000000000000001001","111111111111111100","000000000000000100","000000000000000110","000000000000000110","111111111111111010","111111111111101010","000000000000001001","111111111111111100","000000000000010010","000000000000011111","111111111111111100","111111111111110101","000000000000000000","111111111111110101","000000000000000000","000000000000010111","111111111111101110","000000000000000100","111111111111110101","000000000000010000","111111111111101001","000000000000100010","111111111111110111","000000000000001011","111111111111111001","000000000000001000","111111111111111111","111111111111110111","000000000000011101","000000000000000100","111111111111110000","000000000000100000","111111111111111111","000000000000010111","000000000000010000","000000000000010100","111111111111111001","000000000000001110","000000000000100000","000000000000000011","000000000000000001","111111111111011111","111111111111111011","111111111111011111","111111111111110101","111111111111000100","111111111111111110","111111111111111001","111111111111110001","000000000000000000","000000000000000111","111111111111111010","000000000000010101","000000000000100011","000000000000010010","000000000000011001","000000000000001001","000000000000000000","000000000000011101","111111111111100101","000000000000000100","000000000000010010","111111111111110101","000000000000010000","000000000000000111","000000000000011001","111111111111111011","000000000000000010","000000000000011001","000000000000011101","111111111111100111","000000000000101100","000000000000010101","000000000000110011","000000000000011101","111111111111110100","000000000000010000","111111111111111000","000000000000000010","111111111111110101","000000000000000011","111111111111111100","111111111111111010","000000000000011001","111111111111110000","000000000000011100","111111111111011100","000000000000001100","000000000000100110","111111111111111111","111111111111111001","111111111111101110","111111111111100111","000000000000000110","000000000000000010","000000000000010101","000000000000100100","000000000000001101","000000000000010111","000000000000000111","111111111111110010","111111111111111001","000000000000000000","000000000000011001","111111111111111000"),
("111111111111001111","111111111111110011","111111111111101011","000000000000000110","111111111110100001","111111111111110111","000000000000001001","000000000000011111","000000000000010011","000000000000000000","111111111111101100","111111111111110111","111111111111111000","111111111111010110","111111111111111001","111111111111110011","000000000000000111","000000000000001010","111111111111111010","000000000000000001","111111111111011100","111111111111100111","111111111111101100","111111111111111000","111111111111101001","000000000000011101","000000000000001011","000000000000011000","000000000000011011","111111111111101110","000000000000010100","000000000000000110","000000000000001111","111111111111111000","000000000000000110","000000000000000101","111111111111111000","000000000000100010","000000000000100101","111111111111101011","111111111111111010","111111111111110001","000000000000001110","111111111111101001","000000000000011101","000000000000000000","111111111111111111","000000000000011010","000000000000000000","000000000000010001","000000000000010110","000000000000011001","000000000000010000","111111111111111101","000000000000000000","111111111111110101","000000000000010011","000000000000000101","000000000000011100","000000000000000010","000000000000001000","000000000000011111","111111111111111100","111111111111111010","111111111111110010","000000000000001100","111111111111001110","000000000000010000","111111111111011010","111111111111111101","000000000000001000","111111111111110010","111111111111110001","000000000000011011","000000000000010111","000000000000000100","111111111111111101","000000000000011111","000000000000011111","000000000000001011","000000000000000011","000000000000010111","111111111111100010","111111111111100100","000000000000000010","111111111111110111","111111111111111101","111111111111110011","111111111111111110","000000000000000010","000000000000010011","000000000000000110","000000000000100000","111111111111111001","000000000000010010","000000000000001001","000000000000110111","000000000000010101","000000000000011001","000000000000000001","111111111111110111","000000000000000100","111111111111100101","000000000000011011","000000000000010000","111111111111111111","000000000000100100","111111111111100101","111111111111110011","111111111111110101","000000000000001001","000000000000010000","111111111111111101","000000000000000011","000000000000000110","111111111111011111","000000000000000100","111111111111111000","000000000000010001","111111111111111000","111111111111111111","000000000000010111","111111111111111100","111111111111110100","111111111111110111","000000000000000011","111111111111111011","111111111111111011"),
("111111111111010011","000000000000001010","111111111111000101","000000000000000111","111111111110011000","111111111111101010","000000000000011000","111111111111101100","000000000000101000","111111111111111101","000000000000001101","111111111111110101","111111111111111010","111111111111010011","000000000000001010","000000000000001010","111111111111110100","000000000000011111","000000000000000110","000000000000011000","111111111111101011","000000000000000000","111111111111110000","111111111111111110","000000000000001111","111111111111111011","111111111110111110","000000000000001011","000000000000001111","111111111111111111","111111111111111011","111111111111111100","000000000000011101","000000000000000010","000000000000000101","000000000000000011","000000000000000000","000000000000010011","000000000000010001","000000000000000000","000000000000010100","111111111111110111","111111111111111101","000000000000000001","000000000000010101","000000000000010000","000000000000000111","000000000000000100","000000000000001111","000000000000001110","111111111111110100","111111111111110101","000000000000011111","000000000000000000","000000000000010101","111111111111111100","000000000000010010","000000000000010001","000000000000001011","111111111111110110","111111111111110001","000000000000001000","000000000000011101","111111111111101111","111111111111110000","000000000000010111","111111111111111011","000000000000000100","111111111111011100","000000000000000000","111111111111110010","000000000000001011","111111111111001011","000000000000001000","111111111111111110","000000000000000111","000000000000001101","000000000000011001","111111111111110110","000000000000000100","111111111111101010","000000000000010001","000000000000000000","111111111111000010","000000000000011101","111111111111011001","000000000000001011","111111111111111011","000000000000000010","000000000000000101","000000000000010000","000000000000000010","000000000000100101","000000000000001001","000000000000001111","000000000000011011","000000000000101101","000000000000001001","000000000000001001","111111111111111010","000000000000000100","111111111111111001","111111111111111010","000000000000100100","000000000000000100","000000000000000111","000000000000011001","111111111111111100","111111111111110100","111111111111111100","111111111111110100","000000000000001111","000000000000001100","000000000000010011","111111111111011111","000000000000000011","000000000000000000","000000000000000000","000000000000000111","000000000000001111","000000000000000000","000000000000011101","111111111111111100","111111111111110100","111111111111010111","000000000000001000","111111111111110110","111111111111111010"),
("111111111111100000","000000000000001000","111111111111001011","000000000000011001","111111111111011011","111111111111111010","111111111111110100","111111111111100111","000000000000011110","000000000000000011","111111111111110010","000000000000000111","111111111111111101","000000000000000001","111111111111111000","000000000000000000","111111111111101101","000000000000011111","000000000000001010","111111111111111001","111111111111001001","000000000000000000","000000000000001010","111111111111101111","000000000000001000","111111111111110110","111111111111000010","000000000000100000","111111111111110110","111111111111111110","111111111111111110","111111111111100111","000000000000001101","000000000000001011","000000000000001110","111111111111111000","111111111111110110","000000000000100000","000000000000010011","111111111111101011","111111111111111101","000000000000010110","111111111111100001","000000000000000010","000000000000011001","000000000000101010","111111111111111000","000000000000001110","000000000000011101","111111111111110110","111111111111111101","000000000000000111","000000000000011001","111111111111110100","000000000000000001","111111111111111010","111111111111110101","000000000000010010","111111111111110000","000000000000000001","111111111111110000","000000000000010101","000000000000011011","000000000000001010","111111111111110101","000000000000000110","111111111111101110","000000000000001001","111111111111010010","000000000000000100","111111111111111011","111111111111111000","111111111111100001","000000000000010000","111111111111111110","111111111111101110","000000000000000000","000000000000101000","000000000000001100","000000000000001000","000000000000001010","000000000000010110","111111111111100011","111111111111001101","111111111111111110","000000000000000011","111111111111110111","111111111111110100","111111111111110110","000000000000000000","000000000000100001","000000000000011111","000000000000011010","000000000000011011","000000000000000001","111111111111111000","000000000000010111","111111111111111101","000000000000100011","111111111111111010","111111111111111011","111111111111110000","111111111111100000","000000000000011011","000000000000001101","000000000000011000","000000000000001001","111111111111101000","111111111111111000","000000000000000010","111111111111110001","000000000000001001","000000000000001110","000000000000011010","111111111111111110","000000000000001100","000000000000000010","000000000000010110","000000000000000110","000000000000001000","000000000000000110","000000000000001001","111111111111111000","111111111111100010","111111111111100001","000000000000011001","111111111111101100","111111111111110110"),
("111111111111101100","000000000000000001","111111111111001011","000000000000011110","000000000000000110","111111111111101110","111111111111110111","111111111111110001","000000000000101001","000000000000001010","111111111111101110","111111111111011101","111111111111101100","111111111111100110","111111111111110111","111111111111101100","111111111111111000","000000000000010110","000000000000000111","000000000000010101","111111111111001100","111111111111111101","111111111111110010","000000000000010000","111111111111101110","000000000000010001","111111111111010001","000000000000010010","000000000000000000","000000000000000100","000000000000001000","111111111111111001","111111111111111101","000000000000000111","111111111111101011","000000000000010000","111111111111111110","000000000000010010","111111111111111000","111111111111100111","000000000000001011","000000000000001001","111111111111111100","111111111111111000","000000000000001001","000000000000101000","111111111111111101","111111111111111100","000000000000000100","000000000000000100","000000000000000000","000000000000010100","000000000000000111","111111111111101000","000000000000000101","000000000000001001","000000000000010010","000000000000011000","000000000000001110","111111111111101011","111111111111101100","000000000000010011","000000000000001111","000000000000010010","000000000000000000","000000000000010001","111111111111101111","111111111111101011","111111111111101100","111111111111101001","000000000000010101","000000000000000001","111111111111101110","000000000000000001","111111111111111011","000000000000000111","000000000000001000","000000000000011010","111111111111110000","000000000000000000","111111111111110011","111111111111111100","111111111111111000","111111111111100011","000000000000010111","111111111111111011","111111111111100010","111111111111111101","111111111111111111","000000000000010110","000000000000100000","111111111111111011","000000000000010000","000000000000010110","111111111111110001","000000000000001111","000000000000001110","111111111111101100","000000000000100010","000000000000000011","000000000000001000","111111111111001110","111111111111110011","000000000000000000","111111111111101110","000000000000010010","000000000000000101","111111111111111001","111111111111111001","000000000000001111","111111111111111001","111111111111110010","000000000000011000","111111111111111011","111111111111101110","000000000000011100","111111111111110000","111111111111111101","111111111111110001","000000000000000001","000000000000000111","111111111111110110","000000000000000001","111111111111101011","000000000000000111","000000000000100000","111111111111110110","111111111111111011"),
("000000000000000001","000000000000000000","111111111111010010","000000000000011101","000000000000101101","111111111111111001","000000000000000000","111111111111011110","000000000000001010","111111111111110010","111111111111111101","111111111111111111","111111111111111110","111111111111101111","111111111111101110","000000000000010101","111111111111101111","000000000000010111","000000000000001111","000000000000001100","111111111111010111","111111111111100111","111111111111101001","000000000000000101","111111111111111010","000000000000001100","111111111111001011","000000000000000000","000000000000000111","000000000000001100","000000000000001100","111111111111100101","000000000000010010","111111111111111100","111111111111111000","000000000000011010","111111111111101011","000000000000100101","111111111111010101","000000000000001010","000000000000000101","000000000000011110","111111111111001011","111111111111101100","000000000000001101","000000000000010001","000000000000000001","111111111111111101","000000000000010101","000000000000000000","111111111111101111","000000000000010001","111111111111111101","111111111111010111","000000000000010001","000000000000001011","111111111111101101","000000000000011011","111111111111101011","111111111111110101","111111111111101010","000000000000001011","000000000000011011","111111111111111001","111111111111100010","111111111111111011","111111111111110000","000000000000000001","000000000000000001","111111111111100011","000000000000000110","000000000000010001","000000000000000010","111111111111101111","000000000000000101","111111111111110111","000000000000000000","000000000000100001","111111111111101011","000000000000000001","111111111111010000","000000000000011001","000000000000000000","111111111111110000","000000000000000000","111111111111101100","111111111111110101","000000000000011001","111111111111110001","000000000000000110","000000000000010110","000000000000001110","000000000000000111","000000000000011001","111111111111100010","111111111111110011","000000000000011001","111111111111111110","000000000000001100","111111111111111110","000000000000000000","111111111111011110","000000000000001111","000000000000010010","111111111111111001","000000000000011010","111111111111111111","000000000000000101","111111111111110000","111111111111101001","111111111111101010","000000000000011000","000000000000011110","000000000000010110","000000000000010101","000000000000101001","111111111111110101","000000000000001000","000000000000000000","000000000000010010","000000000000010100","111111111111110001","000000000000000000","111111111111110101","111111111111110011","000000000000011111","111111111111110100","000000000000000001"),
("000000000000001001","000000000000001000","111111111111100001","000000000000011001","000000000000111011","000000000000010010","000000000000000110","111111111111110010","000000000000001001","111111111111101111","111111111111111001","111111111111111111","000000000000000101","111111111111010010","111111111111110001","000000000000001010","000000000000001010","000000000000100001","111111111111110111","111111111111110000","111111111110111101","111111111111110001","000000000000000100","000000000000010101","111111111111101101","000000000000001010","111111111111111001","000000000000000101","111111111111110001","000000000000001100","000000000000000000","111111111111111000","000000000000100011","000000000000011010","111111111111110101","000000000000010001","111111111111101100","000000000000001110","111111111111110010","111111111111111101","000000000000010001","000000000000000111","111111111110111010","111111111111011011","000000000000100110","111111111111100001","000000000000000011","000000000000000100","000000000000010101","111111111111110110","111111111111101011","000000000000001110","000000000000010111","111111111111100001","000000000000001101","000000000000000100","111111111111110000","111111111111111101","111111111111110100","111111111111111010","000000000000000000","000000000000000000","000000000000011111","000000000000000000","111111111111110101","000000000000011100","000000000000001000","111111111111111100","000000000000000010","111111111111110001","111111111111101110","000000000000000000","111111111111010111","111111111111001100","000000000000000111","111111111111101011","000000000000001111","000000000000010101","111111111111110110","000000000000001101","111111111111100001","000000000000000001","000000000000001010","111111111111111010","000000000000001011","111111111111100100","000000000000011100","000000000000000000","000000000000000001","111111111111101100","111111111111101010","000000000000000110","111111111111110001","111111111111111011","111111111111100101","000000000000000101","111111111111111010","111111111111110101","111111111111110001","111111111111100111","000000000000011001","111111111111110111","000000000000001111","000000000000000001","111111111111111001","111111111111111111","111111111111110100","111111111111100011","111111111111111111","000000000000001111","000000000000001100","111111111111111101","000000000000011101","000000000000000000","111111111111110101","000000000000100111","000000000000001100","000000000000000011","000000000000000000","000000000000000001","000000000000000101","000000000000001010","000000000000000001","000000000000010001","111111111111011001","000000000000011101","111111111111111010","111111111111111101"),
("000000000000010101","000000000000000000","111111111111100100","000000000000100100","000000000000100110","111111111111111011","000000000000000000","111111111111100110","111111111111110011","000000000000011001","000000000000010111","111111111111110110","000000000000010101","111111111111101011","111111111111010010","000000000000000011","000000000000100011","000000000000100011","000000000000010000","000000000000011101","111111111111000000","000000000000000001","000000000000100010","000000000000001001","111111111111101100","000000000000000010","000000000000000101","111111111111111000","111111111111110110","000000000000000011","000000000000010011","111111111111101000","000000000000100111","000000000000011110","000000000000000001","111111111111110110","111111111111101100","111111111111101111","111111111111011111","000000000000000000","000000000000000111","000000000000010001","111111111111000011","000000000000000000","111111111111111111","111111111111100111","111111111111011100","111111111111110110","000000000000010011","000000000000001110","111111111111100110","000000000000010000","111111111111110010","000000000000001100","000000000000001010","111111111111111001","111111111111101011","000000000000000001","000000000000010111","000000000000001011","111111111111111000","000000000000001000","000000000000100111","000000000000001010","111111111111110110","111111111111111100","111111111111110001","000000000000011100","111111111111110111","111111111111011111","000000000000010110","111111111111111001","111111111111100010","111111111111010101","000000000000011000","111111111111110011","000000000000010100","000000000000100011","111111111111111111","111111111111111110","111111111111111000","111111111111111001","000000000000001010","111111111111110000","000000000000100111","000000000000010010","000000000000011101","000000000000000000","111111111111101110","000000000000000001","111111111111111100","000000000000011011","111111111111110011","000000000000001101","111111111111101101","000000000000001110","111111111111100010","000000000000000011","000000000000001100","111111111111110100","000000000000000101","111111111111111101","000000000000110001","000000000000000010","111111111111111000","000000000000010011","111111111111111111","111111111111101001","111111111111111011","000000000000001001","111111111111101001","000000000000001111","111111111111111001","000000000000010010","000000000000000100","000000000000011011","000000000000011000","111111111111110100","111111111111101111","000000000000001100","000000000000001001","111111111111111001","111111111111110100","000000000000010001","111111111111110011","000000000000101100","000000000000011011","111111111111111010"),
("000000000000100011","000000000000001000","111111111111011010","000000000000011111","000000000000110000","000000000000000001","111111111111110011","111111111111101001","111111111111110011","111111111111111010","000000000000001010","111111111111110011","000000000000011110","111111111111001100","111111111111011000","000000000000000000","000000000000011100","000000000000000001","000000000000010001","000000000000010011","111111111111001000","111111111111110101","000000000000111111","000000000000000001","000000000000000000","000000000000001011","000000000000010110","111111111111111000","000000000000011100","000000000000000001","000000000000001111","111111111111101010","000000000000001011","000000000000010110","111111111111101111","000000000000100110","111111111111110000","000000000000010000","111111111111010000","111111111111110111","000000000000000011","000000000000000011","111111111111010001","111111111111101111","000000000000000110","111111111111110111","000000000000000011","111111111111111010","000000000000010010","000000000000001101","111111111111111001","111111111111111110","111111111111101011","111111111111111011","000000000000001001","111111111111111111","111111111111111100","000000000000001001","000000000000000000","000000000000001001","000000000000010100","000000000000001000","111111111111111100","000000000000100000","111111111111110001","111111111111110110","111111111111110010","000000000000010111","111111111111111101","111111111111101101","000000000000011100","111111111111110101","111111111111011101","111111111111000110","000000000000011000","000000000000010010","000000000000001011","111111111111110011","111111111111111110","111111111111101110","111111111111110011","111111111111101101","000000000000000110","111111111111110110","000000000000010101","111111111111100010","111111111111111001","111111111111111010","000000000000010011","111111111111011011","111111111111011111","000000000000100100","111111111111011111","111111111111101001","111111111111000100","111111111111110110","111111111111101101","111111111111101101","000000000000000110","111111111111111111","000000000000001011","000000000000000010","000000000000111000","000000000000001110","111111111111111100","000000000000001011","111111111111110011","111111111111101000","111111111111110101","111111111111110110","111111111111101110","000000000000010110","000000000000011111","000000000000001011","000000000000001010","000000000000010001","000000000000001110","000000000000000001","111111111111100011","111111111111110011","111111111111111110","000000000000000000","111111111111100011","000000000000001010","111111111111011010","000000000000101010","111111111111111001","000000000000000001"),
("000000000000011011","111111111111111000","111111111111111011","111111111111111101","000000000000011111","000000000000011101","000000000000000001","111111111111110100","111111111111111011","000000000000000000","111111111111101111","111111111111100111","000000000000001001","111111111111110011","111111111111100100","000000000000100011","000000000000011010","000000000000010111","000000000000010111","111111111111101111","111111111111100000","111111111111100110","000000000000011100","111111111111111110","000000000000000101","000000000000011110","111111111111111010","111111111111100011","000000000000010101","000000000000001001","000000000000010111","111111111111110100","000000000000010010","000000000000100101","111111111111111101","000000000000010111","111111111111110010","000000000000000101","111111111111101100","000000000000000100","000000000000000010","000000000000100101","111111111111101110","000000000000000000","000000000000011110","111111111111010110","111111111111011110","111111111111111111","000000000000001111","111111111111110011","000000000000000111","000000000000010101","111111111111010100","111111111111110100","111111111111101111","111111111111111011","000000000000000101","111111111111110100","111111111111110101","000000000000000100","000000000000000000","000000000000010001","111111111111110101","111111111111111011","111111111111100111","000000000000001110","111111111111111111","000000000000011000","000000000000010011","000000000000001011","000000000000000010","111111111111111001","111111111111111010","111111111110110110","000000000000000101","111111111111110000","000000000000010001","000000000000010001","111111111111101000","111111111111101111","000000000000100011","000000000000011001","111111111111111100","111111111111110010","000000000000100111","111111111111100111","000000000000000000","000000000000011100","000000000000010000","111111111110111101","111111111111100010","000000000000010101","111111111110110110","111111111111101001","111111111111010001","000000000000000101","111111111111000111","000000000000001110","111111111111111010","111111111111111000","111111111111111001","000000000000010111","000000000000100110","000000000000110000","000000000000001101","000000000000000101","000000000000000000","111111111111010011","111111111111100110","111111111111110111","000000000000000101","000000000000010010","000000000000100001","111111111111111110","000000000000010000","000000000000010001","000000000000010011","111111111111111111","111111111111100111","000000000000001000","000000000000001100","111111111111110000","111111111111010011","000000000000000111","111111111111101011","000000000000000001","000000000000001110","111111111111101011"),
("111111111111110111","000000000000011001","111111111111111011","000000000000001011","000000000000011010","000000000000011000","111111111111101101","000000000000011101","111111111111010110","111111111111111110","000000000000010101","000000000000000000","000000000000001001","111111111111110101","111111111111010100","000000000000011101","000000000000001011","000000000000100001","000000000000010111","111111111111110100","111111111111011001","000000000000011001","000000000000010110","111111111111111000","111111111111110101","111111111111111011","000000000000100111","111111111111101110","111111111111101000","111111111111111111","000000000000010110","111111111111011100","111111111111111100","000000000000011011","000000000000000001","000000000000011000","000000000000000001","000000000000001010","111111111111110011","111111111111110011","111111111111111101","000000000000000011","000000000000000001","111111111111110111","000000000000010110","111111111111101011","111111111111101011","111111111111110011","000000000000000111","000000000000001000","000000000000010101","000000000000011010","111111111111101101","000000000000000101","111111111111111101","000000000000010111","111111111111110110","111111111111110011","111111111111011111","000000000000000101","000000000000001010","111111111111111001","000000000000000000","000000000000010001","111111111111001010","111111111111110101","111111111111111011","000000000000011100","000000000000001000","000000000000000000","000000000000001000","000000000000010111","111111111111110001","111111111111000110","000000000000011011","111111111111011001","000000000000010001","000000000000010000","111111111111101111","000000000000000110","111111111111111011","111111111111100100","111111111111110011","111111111111111101","000000000000100000","111111111111100010","111111111111110011","111111111111110010","000000000000000110","111111111111011111","111111111111110011","000000000000000101","111111111110101111","111111111111011000","111111111111101001","111111111111111001","111111111111000011","111111111111110010","111111111111111100","000000000000011011","111111111111110100","000000000000010010","111111111111111110","000000000000101011","000000000000000100","000000000000100110","111111111111111100","111111111111001010","111111111111110011","000000000000001111","111111111111101011","000000000000000110","000000000000100101","111111111111011110","000000000000011110","000000000000000111","111111111111110000","000000000000010001","111111111111101011","111111111111110101","000000000000010010","111111111111111110","111111111111000111","000000000000000010","111111111111100000","111111111111111110","000000000000000010","000000000000000000"),
("000000000000001001","000000000000000001","000000000000010010","111111111111101101","000000000000001110","111111111111111001","111111111111010001","000000000000100000","111111111111010001","000000000000001001","000000000000011000","000000000000010101","111111111111111010","111111111111110111","111111111111011001","000000000000100011","000000000000011011","000000000000000111","111111111111111110","111111111111111011","111111111111100001","000000000000001000","000000000000101010","000000000000000101","000000000000000010","000000000000000001","000000000000100100","111111111111110101","111111111111100011","000000000000010101","000000000000010000","111111111111110100","111111111111110010","111111111111110111","000000000000000111","000000000000000000","111111111111110001","000000000000000000","111111111111110110","000000000000001110","000000000000000000","000000000000010010","111111111111101101","111111111111101111","000000000000010100","111111111111101001","111111111111110100","111111111111101101","000000000000001111","000000000000001100","000000000000101001","000000000000000101","111111111111101001","000000000000000010","000000000000001001","000000000000001010","000000000000000001","000000000000001110","111111111111100101","111111111111111110","111111111111111000","000000000000010111","111111111111101101","000000000000001000","111111111110111101","000000000000000010","111111111111110101","000000000000000011","000000000000000000","111111111111101000","000000000000000000","000000000000000001","111111111111100100","111111111111011101","000000000000000000","111111111111110001","111111111111110100","000000000000011000","111111111111101000","111111111111111011","000000000000010001","111111111111110011","111111111111110001","000000000000010011","000000000000011111","111111111111111010","000000000000011101","000000000000001011","111111111111101100","111111111111110100","111111111111110100","111111111111101101","111111111110111111","111111111111111111","111111111111101101","111111111111110001","111111111110110100","111111111111100100","111111111111110111","000000000000000001","000000000000000010","000000000000011011","000000000000011111","000000000000010111","111111111111100110","000000000000011001","111111111111100110","111111111111010111","000000000000000000","000000000000000100","111111111111100000","000000000000100101","000000000000001110","111111111111100011","000000000000101001","111111111111101110","111111111111111110","000000000000000101","111111111111111111","000000000000000010","000000000000010001","000000000000000011","111111111111100101","111111111111101001","111111111111101100","111111111111110011","000000000000001111","111111111111110011"),
("000000000000010100","111111111111100110","000000000000000101","111111111111011111","000000000000001001","000000000000100100","111111111111010000","000000000000101111","111111111111101011","000000000000000100","000000000000010001","000000000000110001","111111111111111101","111111111111100100","111111111111100010","000000000000001110","000000000000100011","111111111111111101","000000000000000000","111111111111100001","111111111110111110","111111111111111000","000000000000001110","111111111111011010","111111111111101000","111111111111101100","000000000000010111","000000000000000010","000000000000001011","000000000000010000","111111111111101110","111111111111111110","111111111111111001","111111111111111111","000000000000001000","000000000000000111","000000000000001010","000000000000000001","000000000000000101","111111111111110101","000000000000011101","000000000000101001","111111111111111110","111111111111110110","000000000000011010","000000000000010110","111111111111110101","000000000000000100","000000000000001010","000000000000010101","111111111111101100","111111111111110100","111111111111010110","111111111111111001","111111111111110100","111111111111110100","111111111111111110","000000000000000001","111111111111100101","000000000000000100","111111111111101010","000000000000010000","111111111111011110","111111111111111010","111111111111101010","000000000000000011","000000000000000001","000000000000001000","000000000000101100","000000000000010100","111111111111110011","000000000000000010","000000000000000001","111111111111101100","111111111111111101","000000000000000111","000000000000001000","111111111111100111","000000000000000101","000000000000001111","000000000000100010","111111111111110010","000000000000000011","111111111111111110","111111111111101101","000000000000001001","000000000000010010","000000000000001001","000000000000001100","111111111111011111","111111111111111110","111111111111111010","111111111110101010","111111111111100011","111111111111111000","111111111111100001","111111111111010100","111111111111110001","000000000000010110","000000000000101101","000000000000001011","000000000000010011","000000000000010001","000000000000001011","111111111111010010","000000000000001011","111111111111011101","111111111111000100","000000000000000001","000000000000001111","111111111111010011","000000000000100110","000000000000011010","111111111111101010","000000000000010001","000000000000000111","000000000000001100","000000000000001101","111111111111101111","000000000000000110","000000000000100001","000000000000001101","111111111111100111","000000000000001000","000000000000000010","111111111111101001","000000000000000011","000000000000000110"),
("000000000000010001","111111111110111101","111111111111111111","111111111111101011","000000000000000011","000000000000011110","111111111111100101","000000000000001010","000000000000000001","111111111111100010","111111111111101101","000000000000110111","000000000000000100","111111111111100100","111111111111110010","111111111111110010","000000000000001110","111111111111111111","000000000000001110","111111111111011101","111111111111000010","000000000000010011","111111111111110000","111111111111100010","000000000000000010","000000000000001010","000000000000001010","111111111111011110","111111111111110100","000000000000000100","000000000000000101","111111111111101111","111111111111100110","000000000000010100","000000000000010000","000000000000000001","000000000000011000","000000000000000000","111111111111111001","111111111111100111","000000000000011001","000000000000011110","000000000000000010","111111111111110010","000000000000010001","000000000000010010","111111111111110101","000000000000000100","000000000000000101","000000000000010100","111111111111010011","111111111111111000","111111111111011111","000000000000011001","111111111111111001","000000000000001001","000000000000010101","111111111111111110","111111111111100000","111111111111101111","111111111111011101","111111111111011001","111111111110100101","000000000000001110","111111111111011110","000000000000011101","111111111111100110","000000000000011011","000000000000101001","111111111111110111","000000000000000000","000000000000000100","111111111111110110","111111111111011111","000000000000001011","111111111111101011","111111111111111110","111111111111110101","111111111111110100","111111111111101111","000000000000100000","111111111111110011","000000000000000010","000000000000001111","111111111111110110","111111111111110110","000000000000110000","000000000000010000","111111111111110110","111111111111111110","111111111111111100","111111111111111011","111111111111011110","111111111111010000","000000000000001010","000000000000000100","111111111111111000","111111111111011000","000000000000010010","000000000000000010","000000000000010100","000000000000110001","111111111111110110","000000000000010011","111111111111011010","111111111111110011","111111111111101110","111111111111011111","111111111111101101","000000000000011100","111111111111011111","111111111111111110","000000000000010010","111111111111111010","000000000000001111","000000000000000011","111111111111110110","111111111111111100","111111111111100011","111111111111100111","000000000000101000","000000000000011111","111111111111110001","111111111111101111","000000000000000101","111111111111011101","111111111111110111","000000000000000010"),
("000000000000010010","111111111111100100","111111111111111110","000000000000000111","111111111111011001","000000000000000111","111111111111110111","000000000000001111","000000000000000111","111111111110111110","111111111111111011","000000000000110010","000000000000011101","111111111111011101","111111111111111110","000000000000010000","111111111111110011","111111111111111011","000000000000010110","111111111111111101","111111111111011101","111111111111111101","111111111111101110","111111111111110011","000000000000000110","000000000000001100","000000000000000001","111111111111101011","000000000000000010","000000000000010010","000000000000001011","111111111111101001","000000000000010100","000000000000000001","000000000000010101","000000000000101100","000000000000011100","000000000000011010","111111111111101101","111111111111111011","000000000000110100","000000000000001100","000000000000010001","111111111111110100","000000000000101010","000000000000000011","000000000000011101","000000000000101010","000000000000010011","000000000000001110","111111111111100000","000000000000100101","000000000000011101","000000000000110100","000000000000100000","000000000000011000","000000000000011000","111111111111111111","111111111111111011","111111111111101011","000000000000001011","111111111111110111","111111111111000101","111111111111110100","111111111111100001","000000000000101101","111111111111111100","111111111111111001","111111111111111111","000000000000001001","000000000000000001","000000000000001001","111111111111100101","111111111111101111","000000000000000110","111111111111100010","000000000000111010","111111111111111111","000000000000000011","000000000000011011","000000000000000101","000000000000100100","111111111111110001","111111111111001101","111111111111101001","111111111111110000","000000000000111001","111111111111111111","111111111111100111","111111111111010011","111111111111110100","000000000000101001","111111111111011110","111111111111001110","000000000000010011","111111111111111101","111111111111101011","000000000000000000","111111111111110110","000000000000101011","000000000000010111","000000000000111000","000000000000001101","000000000000000001","111111111111110100","000000000000010111","000000000000001100","111111111111111110","111111111111101010","000000000000000010","111111111111111100","111111111111101001","000000000000101110","000000000000010010","000000000000000110","111111111111010111","000000000000011010","000000000001000011","000000000000001111","000000000000101010","000000000000100111","000000000000010000","111111111111111010","111111111111101011","111111111111100100","111111111111101100","000000000000100010","111111111111110101"),
("000000000000100101","111111111111111110","111111111111111111","111111111111011101","000000000000000001","111111111111111101","111111111111111111","000000000000010110","111111111111111010","111111111111101100","111111111111110100","000000000000100101","111111111111111101","111111111111111010","111111111111011101","000000000000001110","111111111111101000","111111111111111111","000000000000001010","111111111111011000","111111111111101001","000000000000000011","111111111111100101","111111111111111110","111111111111111110","000000000000001011","111111111111111001","111111111111101100","000000000000100000","000000000000100011","111111111111110001","111111111111101101","000000000000011000","000000000000010011","111111111111110110","111111111111110100","000000000000010110","111111111111111010","111111111111100101","000000000000000001","000000000000100101","000000000000111011","000000000000011011","000000000000000100","000000000000011001","111111111111100110","000000000000101100","000000000000001011","000000000000000101","000000000000001010","111111111111011001","111111111111110000","111111111111111111","000000000000000000","111111111111101011","000000000000000100","000000000000101000","111111111111100010","111111111111101111","111111111111111010","000000000000100010","111111111111011011","111111111111011010","111111111111111100","111111111111101101","000000000000100111","111111111111110011","000000000000100100","111111111111110110","000000000000001101","111111111111110111","000000000000000011","000000000000100000","111111111111111001","000000000000011011","000000000000001000","000000000000100001","000000000000000000","000000000000000000","000000000000000000","000000000000000000","000000000000101001","111111111111110001","111111111111010101","111111111111101100","111111111111100011","000000000000011110","111111111111110111","111111111111100001","111111111111100001","111111111111101100","000000000000001001","000000000000000100","111111111111011010","000000000000001000","000000000000000011","111111111111101000","000000000000001000","000000000000100001","000000000000001011","000000000000011001","000000000000110110","000000000000000000","111111111111101110","111111111111111000","000000000000010100","000000000000000111","000000000000001100","111111111111010110","111111111111110010","000000000000000011","111111111111100011","000000000000001110","000000000000010100","111111111111110001","000000000000010010","000000000000101100","000000000000100000","111111111111101110","000000000000101110","000000000000000100","111111111111101111","111111111111111001","111111111111110110","111111111111101111","000000000000010110","000000000000011000","111111111111111011"),
("000000000000011001","111111111111110010","000000000000001011","111111111111110100","000000000000010000","000000000000011111","000000000000100010","000000000000000011","111111111111110000","111111111111111101","111111111111111001","000000000000000100","111111111111110100","111111111111011110","000000000000000000","111111111111110010","000000000000001000","111111111111011010","111111111111101110","111111111111011001","111111111111011101","111111111111110110","111111111111111011","111111111111110110","111111111111101100","000000000000001011","111111111111101101","111111111111110010","000000000000010011","000000000000100011","111111111111101001","111111111111101111","000000000000000001","000000000000010011","111111111111011111","000000000000001110","000000000000010011","111111111111110110","111111111111111110","000000000000010100","000000000000010111","111111111111111111","000000000000011101","000000000000001001","000000000000100110","000000000000000001","000000000000011111","000000000000000000","111111111111111001","000000000000011111","111111111111100001","111111111111110100","111111111111111101","000000000000010010","111111111111100011","111111111111101001","000000000000010011","111111111111100110","111111111111101110","111111111111110001","111111111111100111","111111111111101101","111111111111100110","000000000000001110","111111111111110001","000000000000010101","000000000000000000","000000000000011001","111111111111111000","000000000000000000","000000000000000100","111111111111100110","000000000000010101","111111111111111110","111111111111110111","000000000000010001","000000000000011001","111111111111111001","000000000000001011","111111111111111001","000000000000000011","000000000000000011","000000000000000011","111111111111111001","111111111111101110","111111111111101010","000000000000010010","000000000000001011","000000000000010101","111111111111101111","111111111111111000","111111111111111101","111111111111110111","111111111111111001","000000000000001111","111111111111100110","111111111111111111","000000000000000100","000000000000000010","000000000000011001","000000000000101010","000000000000100111","000000000000010100","111111111111011101","111111111111011100","111111111111110110","000000000000001001","000000000000010110","111111111111111110","000000000000100100","111111111111101000","111111111111101111","000000000000001110","000000000000000011","111111111111011110","000000000000000000","000000000000000101","000000000000000111","111111111111110001","000000000000001010","000000000000010110","000000000000000001","000000000000010101","000000000000010000","000000000000001010","000000000000000100","000000000000100000","111111111111111010"),
("111111111111110010","000000000000000111","111111111111110011","111111111111110110","111111111111110100","000000000000000101","000000000000000011","000000000000000000","111111111111110100","000000000000010001","111111111111110110","111111111111110110","111111111111110011","111111111111111001","000000000000000110","000000000000001011","000000000000001110","111111111111111000","000000000000001000","000000000000001000","111111111111110110","000000000000001001","111111111111111110","000000000000000111","111111111111101110","111111111111110011","111111111111111111","111111111111110010","000000000000010100","000000000000001110","000000000000001000","111111111111111011","000000000000001111","111111111111111001","111111111111101110","000000000000010100","000000000000001111","111111111111101111","000000000000010010","000000000000000110","000000000000000000","111111111111111011","111111111111111111","111111111111111000","000000000000000010","000000000000010010","111111111111110011","000000000000000011","111111111111110101","111111111111111111","000000000000001010","000000000000001010","111111111111111111","111111111111111011","000000000000001101","000000000000001110","111111111111111100","111111111111110010","111111111111110010","000000000000010100","111111111111110011","111111111111110001","000000000000000100","111111111111101101","111111111111101111","000000000000000111","111111111111111010","000000000000010000","000000000000000001","000000000000010010","111111111111111111","000000000000000011","111111111111110000","111111111111111001","000000000000000000","000000000000010011","000000000000010001","000000000000000001","000000000000001000","111111111111110011","000000000000000000","000000000000001100","111111111111110111","111111111111111111","111111111111101100","000000000000000000","111111111111101110","111111111111110101","111111111111111111","111111111111101110","000000000000010000","000000000000001010","111111111111111001","111111111111101111","000000000000000000","111111111111110111","000000000000001110","111111111111110001","000000000000010011","111111111111110101","000000000000010100","111111111111110011","000000000000010010","000000000000000000","111111111111110000","000000000000001111","111111111111110011","000000000000000110","000000000000000000","000000000000001110","111111111111111001","000000000000001000","000000000000001110","000000000000010100","111111111111110010","111111111111101110","111111111111101111","000000000000001000","111111111111110101","111111111111111110","000000000000001100","111111111111111000","111111111111110001","000000000000000001","111111111111101100","000000000000000000","000000000000000110","000000000000001101"),
("000000000000000011","000000000000001100","000000000000000000","111111111111111011","111111111111111100","111111111111111100","000000000000000101","111111111111111110","000000000000001100","000000000000000100","000000000000000000","111111111111110100","000000000000000011","111111111111101011","111111111111111100","111111111111111101","000000000000000101","000000000000001011","000000000000010101","111111111111111101","111111111111100011","000000000000010100","000000000000010000","111111111111111000","111111111111100000","000000000000000100","111111111111111000","000000000000000101","000000000000100011","000000000000100010","111111111111110011","000000000000001111","000000000000001010","111111111111111110","000000000000000010","000000000000011101","111111111111101000","000000000000010001","000000000000001000","000000000000010011","000000000000011110","000000000000001001","111111111111110111","111111111111111111","111111111111111101","000000000000001000","000000000000011110","111111111111110110","000000000000000010","000000000000001100","000000000000010011","000000000000000010","111111111111111011","111111111111100101","000000000000011101","111111111111110110","000000000000000111","000000000000010100","111111111111110001","111111111111111010","000000000000001111","000000000000100010","111111111111111110","111111111111110110","000000000000000000","000000000000000011","111111111111110111","000000000000010010","000000000000000100","111111111111101111","111111111111111101","000000000000000011","000000000000011000","000000000000000101","000000000000011110","111111111111111111","111111111111101000","000000000000000011","111111111111110000","111111111111111111","000000000000000000","111111111111111110","111111111111110110","000000000000011010","000000000000011111","111111111111111110","111111111111110101","000000000000100000","111111111111111110","000000000000000011","000000000000001101","000000000000000010","111111111111111111","111111111111111000","111111111111100100","000000000000000001","111111111111111011","000000000000000000","000000000000000001","000000000000011011","111111111111111000","000000000000001000","000000000000000000","000000000000001100","000000000000001011","000000000000001101","111111111111100110","000000000000000110","000000000000010011","111111111111101100","111111111111100010","000000000000000111","000000000000010111","000000000000010101","000000000000001101","000000000000000111","111111111111111010","000000000000000010","111111111111101001","000000000000001111","000000000000000100","000000000000001010","111111111111111010","111111111111101100","000000000000000110","111111111111101010","111111111111101110","000000000000001001"),
("000000000000001010","111111111111101111","000000000000011011","111111111111111001","111111111111110001","111111111111010010","111111111111111001","000000000000000110","000000000000001001","000000000000010111","111111111111101111","000000000000011111","000000000000000111","000000000000000011","111111111111110100","111111111111110100","000000000000000101","111111111111110001","000000000000000010","000000000000001100","000000000000000111","000000000000001000","111111111111100001","111111111111110111","000000000000001011","111111111111110110","000000000000000001","111111111111111111","000000000000000000","000000000000010001","111111111111100010","111111111111111001","000000000000010101","111111111111100001","111111111111111000","000000000000000110","000000000000001100","111111111111110111","000000000000010001","000000000000100110","000000000000001111","000000000000000000","000000000000000111","111111111111101110","111111111111111010","000000000000010110","111111111111111110","111111111111101100","000000000000010100","000000000000100001","000000000000001101","000000000000001110","000000000000010001","111111111111111110","000000000000000111","000000000000000100","111111111111111010","111111111111111011","000000000000011100","111111111111111111","111111111111101101","000000000000001000","000000000000000100","111111111111110101","111111111111101101","000000000000100000","000000000000010100","000000000000010100","000000000000011101","000000000000010100","000000000000000101","000000000000000101","000000000000010010","000000000000011110","111111111111111100","111111111111111001","111111111111101001","000000000000000111","000000000000001111","000000000000001110","111111111111101011","111111111111110011","000000000000000011","000000000000110010","111111111111111111","111111111111111110","000000000000100001","000000000000001011","000000000000011000","000000000000001010","111111111111111101","111111111111110010","000000000000100111","111111111111101101","000000000000000110","111111111111101100","000000000000010001","000000000000010001","000000000000000100","000000000000100111","000000000000000010","000000000000000000","000000000000000111","000000000000000110","000000000000001001","111111111111010111","111111111111110101","000000000000010101","000000000000000000","000000000000100000","111111111111101100","111111111111101100","111111111111111101","000000000000100001","000000000000100000","111111111111111011","111111111111101011","000000000000001101","111111111111101111","000000000000001110","000000000000011101","111111111111110101","111111111111110000","000000000000011001","000000000000000000","000000000000010001","111111111111101110","000000000000000000"),
("000000000000000000","000000000000000001","111111111111110010","111111111111101001","111111111111111011","111111111111110110","111111111111110100","000000000000000111","000000000000001110","000000000000001111","000000000000011000","111111111111101000","000000000000100001","000000000000010111","111111111111111100","111111111111100111","000000000000010110","000000000000000011","000000000000011111","000000000000011110","000000000000011001","000000000000110000","111111111111111111","000000000000011100","000000000000000000","111111111111111001","111111111111100010","111111111111101011","000000000000011101","000000000000010010","111111111111111101","000000000000000001","000000000000001010","111111111111010110","111111111111100110","000000000000001010","000000000000001101","111111111111111110","111111111111101010","000000000000000110","111111111111101101","111111111111010111","000000000000000000","000000000000000000","000000000000001000","111111111111111100","000000000000011010","111111111111110100","111111111111101110","111111111111110100","000000000000010111","111111111111100010","111111111111111101","111111111111111100","000000000000011001","000000000000001101","111111111111110111","000000000000010001","000000000000001110","111111111111110010","000000000000001011","000000000000100000","000000000000010001","000000000000001000","111111111111010101","111111111111111110","000000000000000111","111111111111111111","000000000000000000","111111111111111101","000000000000000101","000000000000000100","000000000000101011","000000000000010000","000000000000000110","000000000000100101","111111111111111100","000000000000010000","000000000000001110","000000000000011001","111111111111110100","111111111111101100","000000000000101010","000000000000010000","000000000000000011","111111111111111101","111111111111110110","000000000000010010","111111111111111010","111111111111111001","111111111111100000","111111111111110111","111111111111110011","000000000000000111","000000000000001101","111111111111110010","000000000000110011","000000000000010111","111111111111110011","000000000000001010","111111111111111110","111111111111100010","000000000000000000","111111111111101010","000000000000000010","111111111111101101","111111111111011101","000000000000001110","000000000000000011","000000000000000010","000000000000000100","111111111111110100","111111111111110101","000000000000000000","111111111111111000","111111111111100111","000000000000000110","000000000000011001","111111111111100100","000000000000000010","000000000000000000","111111111111110110","111111111111011010","000000000000100111","000000000000010000","111111111111101111","111111111111110100","111111111111101010"),
("111111111111100111","000000000000011001","111111111111101000","111111111111100101","111111111111110000","000000000000101010","000000000000010110","000000000000010001","000000000000001000","000000000000010001","000000000000100000","111111111111101001","000000000000000111","111111111111111110","000000000000010000","111111111111101101","000000000000011111","000000000000000111","000000000000001110","000000000000010000","000000000000000000","000000000000011100","000000000000001001","000000000000000110","000000000000001001","000000000000000000","111111111111110011","000000000000001010","000000000000100110","000000000000000011","111111111111101000","111111111111110111","000000000000010000","111111111111001011","111111111111111100","111111111111101110","111111111111111101","111111111111111101","000000000000001011","000000000000011001","000000000000000010","111111111111010000","000000000000000011","111111111111110111","000000000000000110","111111111111111001","000000000000101001","111111111111110000","111111111111101111","000000000000000010","000000000000000000","111111111111111111","111111111111110100","000000000000001101","000000000000001000","111111111111111101","111111111111100101","000000000000011001","111111111111101011","000000000000010011","111111111111110111","111111111111111011","000000000000000100","000000000000000011","111111111111011010","000000000000000000","000000000000100010","111111111111110100","111111111111111101","111111111111110110","111111111111110110","111111111111111100","000000000000110000","111111111111110100","000000000000100000","000000000000001111","111111111111101000","111111111111111011","000000000000000011","000000000000011000","000000000000000000","111111111111011000","000000000000101111","111111111111111100","000000000000000000","000000000000000011","000000000000010110","000000000000011100","000000000000001101","000000000000001111","111111111111101000","111111111111111110","000000000000000110","111111111111100110","000000000000000010","111111111111111110","000000000000011010","000000000000100011","111111111111010001","000000000000000000","000000000000001000","111111111111100010","111111111111101011","111111111111101110","111111111111101110","111111111111101110","111111111111100110","000000000000101101","111111111111110101","111111111111110111","111111111111111111","111111111111101111","000000000000001001","000000000000011000","111111111111010011","111111111111110100","000000000000000101","000000000000011010","111111111111100110","000000000000011110","111111111111110111","000000000000000000","111111111111100110","000000000000010100","000000000000100110","111111111111011101","000000000000000010","111111111111111001"),
("111111111111010001","000000000000001101","000000000000001000","111111111111110100","000000000001000000","000000000000001000","111111111111111101","000000000000000101","111111111111110110","000000000000010011","000000000000000111","000000000000010000","000000000000001000","111111111111100101","000000000000010000","111111111111111010","111111111111111111","000000000000000100","000000000000110100","000000000000000100","111111111111100100","000000000000000001","000000000000000000","000000000000000100","111111111111111000","111111111111110010","000000000000101001","111111111111110001","000000000000010000","111111111111011110","111111111111010110","111111111111110110","000000000000001101","111111111111100000","111111111111110010","111111111111101110","000000000000101100","000000000000010000","000000000000001110","000000000000010001","000000000000110000","111111111111001010","000000000000000111","111111111111110000","000000000000000001","000000000000000000","000000000000010011","111111111111010100","000000000000101011","000000000000010101","000000000000001111","000000000000010001","111111111111111010","111111111111110010","000000000000000000","000000000000001110","111111111111101101","111111111111111100","000000000000001000","000000000000000110","000000000000001100","000000000000011001","000000000000010001","111111111111011101","111111111111110001","111111111111111110","000000000000101101","111111111111011010","000000000000000010","000000000000000010","111111111111010000","000000000000001011","000000000000010001","111111111111111010","111111111111111110","000000000000010111","111111111111100000","111111111111110010","000000000000001011","000000000000000001","000000000000000000","111111111111010011","000000000000100001","111111111111100011","000000000000000101","111111111111111110","000000000000100111","000000000000011011","000000000000000011","000000000000010101","111111111111110110","111111111111101110","000000000000000101","111111111111101010","111111111111011011","111111111111110010","000000000000010101","000000000000000111","111111111111101001","000000000000000111","111111111111011101","111111111111100111","111111111111011111","111111111111101001","000000000000010100","111111111111101001","111111111111111111","000000000000001100","000000000000001100","000000000000100010","111111111111100100","111111111111111010","111111111111110010","000000000000100111","111111111111100101","111111111111101000","111111111111111110","000000000000001010","111111111111100101","000000000000011110","000000000000010101","111111111111111110","111111111111011001","000000000000101000","000000000000101010","111111111111101011","000000000000000100","111111111111110110"),
("111111111111011000","000000000000001010","111111111111011110","111111111111101101","000000000000111011","111111111111011100","000000000000001011","000000000000000010","000000000000011101","000000000000011100","111111111111100000","000000000000001010","000000000000010101","111111111111111100","000000000000101001","111111111111111010","111111111111101101","000000000000011000","000000000000101000","000000000000011000","111111111111111011","111111111111011010","000000000000000101","000000000000001101","111111111111100010","111111111111101011","000000000000010100","111111111111111101","000000000000001000","111111111111011111","111111111111100101","111111111111101111","000000000000001011","111111111110110100","111111111111111001","111111111111111111","000000000000001101","000000000000011001","111111111111100101","000000000000001101","000000000000010011","111111111111101111","000000000000011000","000000000000000111","000000000000000000","111111111111101110","000000000000000010","111111111111011110","000000000000100100","111111111111101111","000000000000010001","111111111111111100","111111111111110111","111111111111110111","000000000000101010","111111111111111011","111111111111011001","000000000000001101","000000000000010000","111111111111101110","000000000000000101","000000000000001001","000000000000011000","111111111111101111","111111111111010001","111111111111110001","000000000000101000","111111111111100110","111111111111111111","111111111111111000","000000000000000000","000000000000110001","000000000000001110","111111111111111110","000000000000000110","111111111111111000","000000000000000000","111111111111100110","000000000000000100","000000000000010011","111111111111111111","111111111111100100","000000000000000000","000000000000010001","000000000000010110","111111111111110010","000000000000000000","000000000000000100","111111111111101111","000000000000010010","111111111111001111","000000000000000110","000000000000000010","111111111111011101","111111111111011110","000000000000000000","000000000000001001","111111111111110111","111111111111011011","000000000000001010","111111111111111110","111111111111111010","111111111111011010","111111111111111011","000000000000000111","111111111111011010","111111111111110111","000000000000011100","000000000000101011","111111111111110111","000000000000001011","000000000000001000","111111111111011110","000000000000010111","111111111111011011","111111111111110110","000000000000001110","000000000000000000","111111111111010001","000000000000010000","000000000000000000","111111111111100110","111111111111110100","000000000000010001","000000000000000111","111111111111010010","000000000000000001","000000000000000000"),
("111111111111001000","111111111111111101","000000000000000000","111111111111101100","000000000000111101","111111111111101011","000000000000001111","000000000000101110","000000000000000011","111111111111111100","000000000000000101","000000000000010011","000000000000001101","111111111111110100","000000000000010110","000000000000000100","111111111111110011","000000000000010100","000000000000010011","111111111111110101","111111111111100000","111111111111011111","000000000000000110","000000000000000011","111111111111011000","000000000000010010","000000000000010001","111111111111111001","000000000000000001","111111111111001001","111111111111010111","111111111111111000","000000000000000000","111111111111011000","000000000000001010","111111111111110110","111111111111111010","111111111111111101","000000000000000010","000000000000001101","000000000000011110","111111111111100101","000000000000001000","111111111111111001","000000000000001100","111111111111101110","111111111111111110","111111111111011000","000000000000000100","111111111111101110","000000000000000000","000000000000001000","000000000000000101","000000000000000001","000000000000000010","000000000000001101","111111111111011000","000000000000010000","000000000000010001","111111111111111001","111111111111111011","000000000000011101","000000000000010110","111111111111011100","111111111111001000","000000000000001000","000000000000000111","111111111111110001","111111111111100101","111111111111110000","111111111111111111","000000000000010101","000000000000000001","111111111111110010","000000000000000000","111111111111110001","111111111111110010","111111111111101111","111111111111111110","111111111111111010","111111111111110110","111111111111111001","000000000000000101","000000000000001101","111111111111101001","111111111111110010","111111111111110110","000000000000000010","111111111111111111","111111111111111100","111111111111011000","000000000000001100","000000000000011101","111111111111110010","111111111111110111","111111111111100101","000000000000010110","000000000000010110","111111111111000000","111111111111110011","111111111111011110","111111111111110101","111111111111101001","000000000000000110","111111111111111001","111111111111100100","111111111111110100","111111111111111100","000000000000010111","111111111111111001","111111111111111010","000000000000010010","000000000000000101","000000000000000000","111111111111011101","111111111111110010","000000000000011000","000000000000001000","111111111111101001","000000000000100000","000000000000000101","111111111111010111","000000000000000110","000000000000001101","111111111111110101","000000000000000100","000000000000010000","000000000000000100"),
("111111111111001001","000000000000000110","111111111111111111","111111111111110110","000000000000111000","111111111111010011","000000000000001001","000000000000000101","111111111111111011","111111111111101010","111111111111111100","000000000000010100","111111111111111010","111111111111110100","000000000000010001","000000000000001111","111111111111100111","000000000000001111","000000000000001101","111111111111111110","111111111111100111","111111111111010111","111111111111100000","111111111111110000","111111111111010110","111111111111111001","000000000000000100","111111111111110100","111111111111111010","111111111111101000","111111111111110100","111111111111101010","111111111111111100","111111111111100010","000000000000000010","000000000000000010","000000000000001010","111111111111101101","000000000000000100","111111111111111101","000000000000000000","111111111111110100","000000000000000100","000000000000000111","000000000000000010","000000000000000101","000000000000000100","111111111111111010","000000000000000101","111111111111111110","000000000000011101","000000000000001010","000000000000001100","111111111111111101","000000000000001101","111111111111111011","111111111111111000","111111111111111100","000000000000000010","111111111111110000","111111111111111101","000000000000010101","000000000000001000","111111111111111000","111111111111010000","000000000000011010","111111111111101110","111111111111110100","000000000000011000","111111111111101001","111111111111101001","000000000000001110","000000000000000110","000000000000000000","000000000000001000","111111111111111010","000000000000001010","000000000000000001","000000000000100011","000000000000000011","111111111111110001","000000000000001010","111111111111100010","000000000000100101","111111111111111001","111111111111111011","000000000000011011","000000000000001000","111111111111110100","111111111111111010","111111111111100010","000000000000000111","000000000000101111","111111111111110001","000000000000011000","111111111111000001","000000000000100011","000000000000101010","111111111111011000","000000000000010010","111111111111100011","000000000000001001","111111111111101101","111111111111100010","111111111111100101","111111111111110110","111111111111111011","000000000000010110","000000000000101011","111111111111111101","000000000000001011","111111111111111111","000000000000001011","111111111111111111","111111111111100111","111111111111011100","000000000000001000","111111111111111011","111111111111011001","000000000000001011","000000000000010011","111111111111110110","111111111111111011","000000000000001110","000000000000010001","000000000000000100","000000000000001101","000000000000000000"),
("111111111110111100","000000000000001110","111111111111101110","000000000000000000","000000000000000100","111111111111101001","111111111111111110","000000000000100111","111111111111111010","111111111111111001","111111111111110000","111111111111111101","000000000000001111","111111111111110010","000000000000011111","000000000000000000","000000000000000000","111111111111110110","000000000000000001","000000000000001111","111111111111011110","111111111111100011","111111111111110111","111111111111011001","111111111111100001","000000000000001000","000000000000101110","000000000000001110","111111111111110101","111111111111111111","111111111111110100","000000000000011000","111111111111111100","111111111111111100","000000000000011000","000000000000001110","000000000000001110","111111111111110001","000000000000000010","111111111111111000","000000000000001000","111111111111110101","111111111111111001","111111111111101100","000000000000001101","000000000000000000","111111111111110101","111111111111110100","000000000000100101","000000000000010011","000000000000000001","000000000000010001","111111111111100011","111111111111111110","000000000000011101","000000000000010100","000000000000001001","000000000000000011","000000000000000011","000000000000001101","000000000000000111","000000000000000110","000000000000000111","111111111111100110","111111111111001011","111111111111111001","111111111111110110","111111111111111000","000000000000000111","111111111111001010","111111111111111100","000000000000011101","000000000000000000","111111111111111001","000000000000010110","000000000000001001","111111111111110111","000000000000011100","000000000000001011","000000000000010111","111111111111010000","000000000000010000","111111111111100100","000000000000101010","000000000000000100","000000000000001100","000000000000011011","000000000000000100","000000000000000100","111111111111111101","111111111111100101","111111111111111010","000000000000011100","111111111111100001","000000000000001111","111111111111101001","000000000000101010","000000000001000011","111111111111110011","111111111111110000","111111111111011000","000000000000000101","111111111111011110","000000000000000001","111111111111110000","111111111111101011","000000000000010100","111111111111110111","000000000000011110","111111111111101101","111111111111110001","000000000000001100","000000000000010010","000000000000011001","111111111111111111","111111111111011000","000000000000000001","111111111111110101","111111111111100011","000000000000100011","000000000000000111","111111111111101100","000000000000100010","000000000000000100","000000000000000010","111111111111111111","000000000000000000","000000000000000000"),
("111111111111010000","000000000000011011","111111111111111011","111111111111101000","111111111111010100","111111111111001100","000000000000001001","000000000000010110","000000000000010110","111111111111111011","000000000000000001","000000000000011001","000000000000001111","111111111111101001","111111111111110111","000000000000100100","111111111111110101","000000000000001111","111111111111111111","000000000000000000","111111111111110000","111111111111100011","111111111111101000","111111111111100000","111111111111101001","000000000000001101","000000000000011110","000000000000010111","000000000000000101","000000000000001110","000000000000000001","000000000000001110","111111111111111101","000000000000001010","000000000000010000","000000000000010011","111111111111111010","111111111111110000","000000000000000100","000000000000000000","000000000000001001","111111111111110100","000000000000000011","111111111111101001","000000000000001100","000000000000000001","111111111111101001","111111111111111111","000000000000011011","000000000000001011","000000000000010010","111111111111110101","000000000000010100","000000000000011101","000000000000001110","000000000000000110","000000000000000000","000000000000010010","111111111111111111","111111111111110001","111111111111101000","000000000000100001","000000000000011100","111111111111110000","111111111110110101","000000000000001100","111111111111100001","111111111111100111","111111111111111011","000000000000000100","111111111111111111","000000000000100011","000000000000001010","000000000000010011","000000000000011110","000000000000000000","111111111111111000","000000000000001011","111111111111111010","000000000000010101","111111111111101001","000000000000010011","111111111111100111","000000000000100101","000000000000010011","111111111111101110","000000000000010000","000000000000011000","111111111111110001","000000000000001001","000000000000001000","000000000000000110","000000000000001100","111111111111011110","111111111111111111","111111111111110100","000000000000011101","000000000000001010","111111111111011001","111111111111110111","111111111111111001","111111111111110011","111111111111011111","111111111111111110","111111111111110101","000000000000000101","000000000000010001","111111111111111110","000000000000011100","111111111111110110","000000000000000011","000000000000100100","111111111111110110","000000000000000101","000000000000000111","111111111111101010","000000000000000001","000000000000000100","000000000000011000","000000000000001110","000000000000011011","111111111111111101","000000000000010000","111111111111111011","111111111111110011","000000000000000010","000000000000010101","000000000000000011"),
("111111111111011010","000000000000001100","111111111111011101","111111111111101111","111111111110011100","111111111111110101","000000000000001110","000000000000010111","000000000000001101","111111111111110100","111111111111101111","000000000000000111","000000000000000011","111111111111111000","000000000000001110","000000000000000000","111111111111110000","000000000000001000","000000000000001101","000000000000011000","000000000000000000","111111111111111100","111111111111101110","000000000000001000","111111111111111100","000000000000010001","111111111111110011","000000000000010111","000000000000000110","000000000000000101","000000000000011011","111111111111111001","000000000000010100","111111111111111110","111111111111101110","111111111111111101","000000000000001100","111111111111100110","000000000000101001","111111111111101110","111111111111110011","111111111111111101","000000000000010011","000000000000000110","111111111111110100","000000000000001101","111111111111101010","000000000000010100","000000000000000010","111111111111110000","000000000000000000","111111111111110000","000000000000011001","000000000000101110","000000000000011001","111111111111101011","000000000000001101","000000000000010001","000000000000011011","111111111111101101","111111111111111101","000000000000011011","000000000000011100","111111111111101001","111111111111001111","000000000000011110","111111111111101101","111111111111101001","111111111111111100","111111111111111101","000000000000001111","000000000000000001","111111111111111011","000000000000000001","000000000000001010","000000000000000000","000000000000010010","000000000000001001","111111111111111101","000000000000001010","111111111111110111","000000000000001110","111111111111110111","000000000000001010","000000000000000001","000000000000000001","000000000000000001","000000000000001010","111111111111100111","000000000000100011","000000000000100101","000000000000011110","000000000000100010","111111111111100101","000000000000011100","111111111111111111","000000000000010001","000000000000001101","000000000000010001","000000000000000000","111111111111101100","000000000000011110","111111111111100001","111111111111111111","000000000000001001","111111111111101001","000000000000001111","000000000000010010","000000000000010010","111111111111111111","111111111111111011","000000000000001100","000000000000000011","000000000000010011","000000000000000111","111111111111001000","111111111111110101","000000000000001111","000000000000001110","000000000000100010","111111111111111011","000000000000010010","000000000000010110","000000000000000001","000000000000000000","000000000000001000","111111111111110101","111111111111111110"),
("111111111111010111","000000000000000011","111111111111101010","111111111111111010","111111111110000110","111111111111110010","000000000000001110","000000000000001101","000000000000011000","000000000000000111","111111111111111000","000000000000011001","000000000000011011","111111111111100100","000000000000010111","000000000000010011","111111111111011101","000000000000010001","000000000000010000","111111111111111001","111111111111100101","111111111111101000","000000000000000010","111111111111110111","111111111111110011","000000000000001000","111111111111110010","000000000000100111","000000000000001010","000000000000001100","000000000000000101","000000000000000100","000000000000001011","000000000000000100","111111111111111101","000000000000010111","000000000000000000","000000000000001010","000000000000011010","111111111111111100","000000000000001110","000000000000001001","000000000000010000","111111111111110111","000000000000000001","000000000000010011","111111111111101000","111111111111111001","000000000000000110","000000000000001101","000000000000100011","000000000000001010","000000000000100010","000000000000010001","111111111111110111","111111111111110110","000000000000010111","000000000000100000","000000000000001000","000000000000000000","111111111111010100","000000000000011100","000000000000101000","111111111111100011","111111111111101011","000000000000010101","111111111111100000","111111111111110001","000000000000000101","000000000000001100","000000000000001110","111111111111110110","111111111111011101","111111111111111010","000000000000010100","111111111111101101","000000000000001011","000000000000011010","000000000000000111","000000000000010000","111111111111100110","000000000000000000","111111111111100110","111111111111101101","000000000000000101","111111111111111110","111111111111111000","111111111111100101","000000000000000100","111111111111111000","000000000000010011","000000000000010110","000000000000001110","111111111111110111","000000000000001111","000000000000001001","000000000000010100","000000000000000111","000000000000000100","000000000000001110","111111111111011111","111111111111110100","111111111111011011","000000000000000000","111111111111111001","111111111111110000","000000000000001010","000000000000000110","000000000000001000","111111111111111100","000000000000000110","000000000000100110","000000000000001100","000000000000010101","000000000000001110","111111111111010000","111111111111110011","111111111111111110","000000000000010111","000000000000010101","000000000000100101","000000000000001001","000000000000100000","111111111111111001","111111111111011111","000000000000011001","000000000000010100","000000000000010110"),
("111111111111011010","111111111111110011","111111111111110100","000000000000000000","111111111110010110","111111111111110001","000000000000001110","000000000000001011","000000000000000111","000000000000000000","111111111111110110","000000000000000101","000000000000001110","111111111111100011","000000000000000100","000000000000001001","111111111111101101","000000000000010100","111111111111100011","000000000000001011","111111111111110000","111111111111110110","111111111111110000","000000000000001011","000000000000000110","000000000000001011","111111111111001000","000000000000100001","111111111111110110","000000000000101101","111111111111111001","000000000000000110","000000000000011011","000000000000000110","111111111111111110","000000000000010011","111111111111111011","000000000000000110","000000000000011011","111111111111101010","111111111111111111","000000000000000001","000000000000010110","000000000000000000","000000000000010000","000000000000000011","111111111111111010","111111111111011100","000000000000001000","111111111111110000","000000000000000000","000000000000000101","000000000000011010","000000000000100111","000000000000000011","000000000000000101","000000000000000011","000000000000001101","000000000000010110","000000000000000101","111111111111100110","000000000000100011","000000000000010001","111111111111100011","000000000000001001","111111111111111100","111111111111111001","111111111111101111","000000000000000010","111111111111111000","111111111111110011","000000000000001011","111111111111001111","000000000000000110","000000000000001000","000000000000011001","111111111111110100","000000000000110010","111111111111110100","111111111111110101","000000000000000100","000000000000000111","111111111111100110","111111111111001010","000000000000010001","111111111111111000","111111111111100110","000000000000000100","111111111111101101","000000000000010010","000000000000010001","000000000000010111","000000000000100001","000000000000000110","000000000000001010","000000000000010000","000000000000100000","000000000000001101","000000000000101011","000000000000001110","111111111111110000","000000000000000000","111111111111101000","000000000000000000","000000000000010001","000000000000000111","111111111111111011","111111111111110111","111111111111101010","000000000000001011","000000000000001100","000000000000000110","111111111111101110","111111111111111001","000000000000000000","111111111111001111","000000000000001100","000000000000000011","111111111111111011","000000000000100110","000000000000000100","000000000000010101","000000000000000111","111111111111100101","111111111111101001","000000000000101110","000000000000001011","000000000000010010"),
("000000000000001000","000000000000001101","000000000000001011","000000000000010111","111111111111001101","111111111111111101","000000000000010110","111111111111110000","111111111111111100","000000000000000110","111111111111111011","111111111111111101","000000000000101000","000000000000000011","111111111111100111","000000000000000101","111111111111011011","000000000000100011","111111111111100110","000000000000011101","111111111111011101","111111111111110100","111111111111100110","000000000000010111","111111111111111011","000000000000001101","111111111110110111","000000000000011111","111111111111110011","000000000000001001","111111111111111100","000000000000001110","000000000000010011","000000000000100101","111111111111101000","000000000000001000","000000000000010100","000000000000011010","111111111111111111","000000000000000101","000000000000000001","111111111111111111","111111111111111110","000000000000011000","000000000000010101","000000000000000101","111111111111101011","111111111111011110","000000000000001000","111111111111111110","000000000000000101","111111111111111010","000000000000000101","000000000000100010","000000000000000000","000000000000010101","000000000000001001","000000000000001101","111111111111111011","111111111111110011","111111111111100011","000000000000101001","000000000000101010","111111111111011011","000000000000010110","000000000000001101","000000000000011001","111111111111101111","000000000000000110","000000000000000000","111111111111101100","000000000000000011","111111111111100001","000000000000011101","000000000000010110","111111111111110110","000000000000000000","000000000000111010","000000000000000110","111111111111111110","000000000000000100","000000000000000000","111111111111100101","111111111111001010","000000000000001100","000000000000000010","111111111111111100","111111111111110000","000000000000000110","000000000000001000","000000000000011000","000000000000011110","000000000000001101","000000000000011101","000000000000000100","000000000000101010","111111111111111001","111111111111111000","000000000000100001","000000000000000101","000000000000000101","111111111111101111","000000000000010000","111111111111110101","111111111111110101","111111111111110101","111111111111111011","111111111111111001","111111111111111111","111111111111111011","000000000000000110","000000000000010101","000000000000010000","000000000000000000","000000000000000000","111111111111100001","000000000000000111","000000000000010100","000000000000001000","000000000000001001","111111111111111010","000000000000000110","111111111111111110","111111111111001100","111111111111011110","000000000000111000","000000000000000011","000000000000001111"),
("000000000000000000","111111111111111010","111111111111110110","000000000000010111","000000000000001010","111111111111111100","000000000000000011","000000000000000100","000000000000010101","111111111111111010","000000000000001001","000000000000000001","000000000000101001","111111111111100000","111111111111111110","111111111111111010","111111111111010101","000000000000001111","000000000000010010","111111111111111001","111111111110111110","111111111111101100","111111111111101111","111111111111111101","111111111111111100","000000000000000111","111111111111010001","000000000000110011","111111111111100011","000000000000000110","000000000000000111","000000000000000011","000000000000011100","000000000000011101","111111111111111010","111111111111110101","000000000000000000","111111111111111111","111111111111010110","111111111111111101","000000000000000110","000000000000011011","000000000000000000","000000000000010001","000000000000001000","000000000000001010","000000000000001101","111111111111101110","000000000000000011","111111111111110000","111111111111111000","111111111111111101","000000000000001101","000000000000011000","000000000000000000","111111111111110011","000000000000001001","000000000000000010","000000000000010001","111111111111110010","000000000000000100","000000000000010100","000000000000100100","000000000000001000","111111111111110111","000000000000000110","000000000000001000","000000000000001010","000000000000011011","111111111111001100","000000000000001001","000000000000001000","111111111111001101","000000000000000101","000000000000000101","000000000000001001","000000000000011010","000000000000110011","111111111111110001","111111111111100101","000000000000000000","111111111111111111","111111111111100111","111111111111100011","111111111111111001","000000000000000100","111111111111111110","000000000000000101","111111111111110100","000000000000010010","000000000000000011","000000000000001000","000000000000000000","000000000000010011","000000000000010001","000000000000011111","111111111111110111","000000000000001110","000000000000001001","000000000000000000","000000000000000110","111111111111010111","000000000000010110","000000000000010011","000000000000000101","111111111111111100","000000000000010010","000000000000001011","111111111111010011","000000000000001000","111111111111101110","000000000000010111","000000000000011001","111111111111111100","111111111111110110","000000000000001010","111111111111111000","111111111111111001","111111111111111110","000000000000011001","000000000000000010","111111111111101011","000000000000001001","111111111111101010","111111111111101111","000000000000101010","000000000000010101","000000000000010001"),
("111111111111111100","111111111111101110","111111111111111100","000000000000011010","000000000000111101","111111111111101000","000000000000000101","111111111111011100","000000000000000010","111111111111111111","111111111111100111","000000000000000000","000000000000100101","111111111111111000","000000000000010001","000000000000010001","111111111111010111","000000000000001101","111111111111111111","000000000000000000","111111111111000001","000000000000000000","000000000000000000","111111111111111010","000000000000000100","000000000000010110","111111111111001001","000000000000111111","111111111111110101","111111111111111101","000000000000001001","000000000000000010","000000000000000111","000000000000011001","111111111111110110","000000000000001000","111111111111110111","111111111111110001","111111111111110000","111111111111110111","000000000000000000","000000000000010100","111111111111111010","000000000000000110","000000000000000000","111111111111111001","111111111111100110","111111111111101101","000000000000001100","111111111111110111","000000000000000011","111111111111111000","111111111111111000","000000000000000000","000000000000011001","000000000000000001","111111111111110011","000000000000000101","000000000000000011","111111111111110011","000000000000000110","000000000000001110","000000000000011001","000000000000000111","000000000000000100","000000000000010011","111111111111101101","000000000000001001","000000000000001001","111111111110111111","000000000000001010","111111111111110010","111111111111110000","000000000000100111","000000000000001110","000000000000000111","000000000000010011","000000000000111010","111111111111110001","111111111111111000","111111111111100111","000000000000011111","111111111111110000","111111111111111101","000000000000001010","111111111111111100","111111111111110110","111111111111110101","111111111111111110","000000000000000011","111111111111100111","000000000000011011","111111111111110000","000000000000010100","000000000000010100","000000000000100010","000000000000010010","111111111111111010","000000000000000111","000000000000001100","111111111111111100","111111111111100101","000000000000100001","111111111111110011","111111111111101100","111111111111101011","000000000000000110","000000000000011101","111111111111101000","111111111111111111","111111111111110010","000000000000001110","000000000000001001","000000000000000000","000000000000000110","000000000000110101","000000000000001101","111111111111101101","111111111111110100","000000000000000001","000000000000000000","111111111111111001","111111111111110010","111111111111110100","000000000000000000","000000000000110010","000000000000000110","000000000000001001"),
("000000000000010110","111111111111011001","000000000000000010","000000000000110000","000000000001000011","000000000000000001","000000000000011111","111111111111001001","111111111111111101","111111111111100011","111111111111110010","111111111111110100","000000000000100010","111111111111110100","111111111111110110","000000000000001011","111111111111100100","000000000000000001","000000000000001001","000000000000000111","111111111111011100","111111111111111010","111111111111111111","000000000000000101","111111111111110001","111111111111111111","111111111111001111","000000000000001011","111111111111110101","000000000000001001","000000000000000001","000000000000000101","000000000000100101","000000000000100101","111111111111100111","111111111111101110","000000000000001100","111111111111110010","111111111111100110","111111111111110111","111111111111110100","000000000000000100","111111111111001111","000000000000001101","000000000000001010","111111111111101100","111111111111110110","111111111111011000","000000000000001000","000000000000011001","000000000000000000","000000000000001001","000000000000000000","000000000000000000","111111111111111010","000000000000000000","000000000000001110","000000000000010110","000000000000100010","111111111111111111","000000000000010011","000000000000011111","000000000000001100","111111111111110101","000000000000011000","000000000000001000","111111111111111101","111111111111100111","000000000000000101","111111111111011010","000000000000010011","111111111111111000","111111111111011100","000000000000010000","111111111111111111","000000000000001010","000000000000001001","000000000000101101","000000000000010011","111111111111100010","111111111111110101","111111111111111101","111111111111100110","000000000000001000","000000000000001101","111111111111101101","111111111111110100","000000000000001001","111111111111101000","111111111111111000","111111111111011111","000000000000010001","111111111111001010","111111111111110110","000000000000000100","000000000000111101","111111111111101110","000000000000010001","111111111111111100","111111111111111100","111111111111110101","000000000000000011","000000000000010001","111111111111110111","111111111111111000","111111111111111010","000000000000010011","000000000000011100","000000000000000110","000000000000001001","000000000000010001","111111111111110011","111111111111111110","111111111111111011","000000000000010000","000000000001000001","000000000000001011","000000000000010011","111111111111100011","000000000000000001","000000000000001000","000000000000010001","000000000000010011","000000000000001101","111111111111100101","000000000000010101","000000000000011000","000000000000001110"),
("000000000000101001","111111111111111011","111111111111101100","000000000000011111","000000000000101000","111111111111110000","000000000000000000","111111111111101001","111111111111111110","000000000000000010","111111111111110000","111111111111111111","111111111111111110","111111111111111010","111111111111111101","000000000000000000","111111111111110111","000000000000011111","111111111111111000","000000000000001101","111111111111110111","000000000000010010","000000000000100001","111111111111111110","000000000000000010","000000000000000000","111111111111111101","000000000000001001","000000000000011001","111111111111111110","000000000000011011","111111111111100101","000000000000000100","000000000000101000","111111111111111011","111111111111110100","000000000000001101","111111111111101110","111111111111100111","000000000000000001","111111111111111011","111111111111101001","111111111110110011","111111111111011111","000000000000001100","111111111111111011","111111111111101011","111111111111011110","000000000000010011","000000000000000110","000000000000001000","111111111111111011","111111111111110001","000000000000000011","000000000000011001","111111111111111111","000000000000001011","000000000000010000","000000000000001000","111111111111110000","000000000000101001","000000000000000111","000000000000000100","000000000000000000","000000000000000101","000000000000000000","111111111111111010","111111111111100100","000000000000000001","111111111111101011","111111111111110111","000000000000011000","111111111111101110","111111111111111000","000000000000001000","000000000000010001","111111111111111110","000000000000110110","111111111111101000","111111111111011011","000000000000000010","000000000000000101","000000000000001011","000000000000000010","000000000000001100","111111111111110001","111111111111111011","000000000000010111","111111111111111000","111111111111110101","111111111111011110","000000000000010101","111111111110101011","000000000000001001","000000000000000000","000000000000011100","111111111111110100","000000000000000001","111111111111111010","111111111111110110","000000000000000011","000000000000000101","000000000000011010","111111111111111011","111111111111111101","000000000000000101","000000000000001000","000000000000000000","000000000000000011","111111111111111011","000000000000001000","111111111111110100","111111111111101001","111111111111101100","000000000000001010","000000000001000100","111111111111110100","000000000000000000","111111111111011001","000000000000000001","000000000000101010","111111111111110110","000000000000000101","000000000000001100","111111111111101001","000000000000010100","000000000000001111","000000000000010010"),
("000000000000101011","000000000000001100","000000000000001101","000000000000011101","000000000000000110","111111111111110001","111111111111111110","000000000000000101","000000000000000010","111111111111100010","000000000000000111","000000000000001110","000000000000001100","111111111111110101","111111111111111001","111111111111110010","000000000000010011","000000000000000100","000000000000001100","111111111111110111","111111111111110010","000000000000010000","000000000000010100","000000000000011001","111111111111111100","000000000000010011","000000000000001010","111111111111110010","000000000000011000","111111111111111100","000000000000010011","111111111111110000","000000000000011010","000000000000010101","000000000000001000","111111111111110110","000000000000010100","111111111111101001","111111111111100011","000000000000010101","111111111111110101","111111111111110100","111111111111000111","111111111111101110","000000000000010101","111111111111101101","111111111111010100","111111111111100101","000000000000000000","000000000000001000","111111111111100101","000000000000010000","000000000000000111","111111111111101011","000000000000000011","000000000000100110","000000000000010001","111111111111110000","000000000000010100","111111111111111001","000000000000110000","000000000000011000","000000000000000100","000000000000001110","111111111111100000","000000000000100001","000000000000000000","111111111111111100","000000000000001100","111111111111111100","000000000000010011","000000000000010100","111111111111111011","111111111111001000","000000000000010001","000000000000000101","000000000000001101","111111111111111011","111111111111110101","111111111111101001","000000000000000010","000000000000001101","000000000000000101","000000000000010000","111111111111111110","111111111111100001","000000000000000001","000000000000011011","111111111111110101","111111111111010101","111111111111011111","000000000000100101","111111111110011100","111111111111010010","111111111111100011","000000000000101010","111111111111010111","111111111111111101","111111111111100111","000000000000010110","111111111111101010","000000000000010011","000000000000100001","000000000000011011","111111111111111011","000000000000000110","111111111111111111","111111111111101100","000000000000000101","111111111111100111","000000000000001110","000000000000001110","111111111111110001","000000000000001001","000000000000000011","000000000000001011","111111111111111000","000000000000010011","111111111111111010","000000000000001011","000000000000011011","000000000000000111","000000000000010000","111111111111111000","111111111111011101","111111111111110111","000000000000000011","000000000000000110"),
("000000000000111100","000000000000001011","000000000000001000","111111111111110100","000000000000010111","111111111111111100","111111111111111001","000000000000010010","111111111111100010","111111111111100100","000000000000001011","111111111111101101","000000000000000010","000000000000001100","111111111111111101","111111111111101110","000000000000001001","000000000000011010","000000000000000011","111111111111111111","111111111111101011","111111111111111100","000000000000110111","000000000000011011","111111111111110101","111111111111111111","111111111111111001","111111111111101100","000000000000010011","111111111111111010","000000000000000001","111111111111011000","111111111111101101","000000000000100110","111111111111101100","000000000000001110","111111111111111100","000000000000000010","111111111111110010","000000000000000111","000000000000000101","000000000000001000","111111111111010001","111111111111111001","111111111111110111","111111111111110010","111111111111111111","111111111111100101","000000000000000000","000000000000000011","111111111111101000","111111111111110100","000000000000000001","111111111111101100","111111111111110000","111111111111111111","000000000000010010","000000000000000010","000000000000000111","111111111111111110","000000000000011110","111111111111110010","111111111111101110","000000000000010010","111111111111011110","111111111111111100","000000000000010100","000000000000000111","000000000000000011","111111111111100111","111111111111110001","111111111111110110","000000000000000110","111111111111001010","111111111111111100","111111111111101101","000000000000011000","000000000000001010","000000000000000100","000000000000000011","000000000000010100","111111111111110000","000000000000000010","000000000000000110","000000000000011010","111111111111100001","111111111111111010","000000000000010101","111111111111111010","111111111111011110","111111111111011001","000000000000000010","111111111110010101","111111111111011111","111111111111110010","000000000000010011","111111111111000101","111111111111110001","111111111111111000","000000000000100110","111111111111110000","111111111111101111","000000000000101010","000000000000011111","000000000000001111","000000000000001001","000000000000001010","000000000000000011","111111111111110101","000000000000001001","111111111111110011","000000000000001101","111111111111110111","111111111111111111","000000000000010101","111111111111111100","111111111111111100","111111111111111111","000000000000001001","111111111111111111","000000000000011101","111111111111101110","111111111111110000","000000000000010100","111111111111011101","000000000000000100","000000000000100000","000000000000000000"),
("000000000000011010","000000000000000000","000000000000010011","111111111111111100","111111111111111000","111111111111110100","111111111111110100","000000000000001010","111111111111110000","111111111111110101","000000000000010000","000000000000001011","000000000000001100","000000000000000101","111111111111110111","111111111111111100","000000000000001001","111111111111111001","000000000000010101","111111111111111010","000000000000001000","000000000000011100","000000000000100000","000000000000011101","000000000000000101","111111111111101000","111111111111111000","111111111111101101","000000000000001000","000000000000000100","111111111111101100","111111111111101100","111111111111101101","000000000000011101","111111111111111000","000000000000001110","000000000000000001","000000000000000000","111111111111110110","111111111111111100","111111111111111111","000000000000001011","111111111111101100","111111111111101110","111111111111101010","111111111111111111","000000000000000001","111111111111011011","111111111111101111","000000000000001000","000000000000001010","111111111111111001","000000000000000001","111111111111011111","111111111111110110","111111111111111001","000000000000000101","000000000000001010","000000000000100010","000000000000000111","000000000000010001","111111111111111011","000000000000000000","000000000000000000","111111111111100011","000000000000010011","111111111111110000","111111111111111010","000000000000001000","111111111111110101","000000000000001000","000000000000001010","111111111111111000","111111111111001100","111111111111101010","111111111111110001","111111111111101101","000000000000010100","000000000000000010","000000000000000100","111111111111110100","111111111111111101","000000000000010111","000000000000000111","000000000000011000","000000000000010000","000000000000010101","000000000000001111","000000000000001111","111111111111000000","111111111111111011","000000000000001110","111111111110010111","111111111111111000","000000000000001001","111111111111111100","111111111111010010","111111111111010010","111111111111101001","000000000000101101","111111111111110111","111111111111110011","000000000000000000","111111111111111110","000000000000001000","000000000000000111","000000000000000000","111111111111101110","111111111111111111","111111111111111010","000000000000001001","000000000000001010","000000000000000100","111111111111110100","111111111111110010","000000000000100101","000000000000000110","000000000000000101","000000000000000000","000000000000001111","000000000000100000","111111111111110011","000000000000001000","000000000000011110","000000000000000110","111111111111100001","000000000000001111","111111111111111101"),
("000000000000010101","111111111111110011","111111111111111111","000000000000000010","111111111111100011","111111111111110101","111111111111111000","000000000000011011","111111111111011110","111111111111111101","111111111111111101","000000000000000001","000000000000001111","000000000000010101","111111111111010101","000000000000001011","000000000000100111","000000000000000110","111111111111110011","000000000000010000","111111111111111101","000000000000101110","000000000000001101","000000000000000110","000000000000011001","111111111111111000","000000000000000011","111111111111001111","111111111111010100","000000000000000011","111111111111110001","111111111111010101","111111111111111110","000000000000011110","111111111111111001","111111111111101110","000000000000001111","111111111111110101","000000000000000000","000000000000010011","000000000000001111","111111111111111110","000000000000000001","111111111111101000","111111111111110111","000000000000001001","111111111111011111","111111111111011110","000000000000010010","000000000000000001","000000000000100101","000000000000001110","111111111111111000","111111111111011101","111111111111110101","000000000000010101","111111111111110101","000000000000010100","111111111111111010","000000000000001001","000000000000010001","000000000000010111","111111111111111011","111111111111110100","111111111111001110","000000000000001011","000000000000001101","000000000000001000","111111111111111101","000000000000001001","111111111111110110","000000000000010001","111111111111110111","111111111111001000","111111111111111100","111111111111100001","000000000000001110","111111111111110110","000000000000000011","000000000000001001","000000000000011110","111111111111101000","000000000000000000","000000000000001111","111111111111110111","111111111111111110","000000000000001111","000000000000000101","111111111111101110","111111111111001110","000000000000000011","111111111111111010","111111111110011101","111111111111101111","111111111111110011","111111111111011110","111111111111001000","111111111111010101","111111111111100000","000000000000001001","111111111111101001","000000000000100000","000000000000000001","000000000000001001","000000000000000011","111111111111111000","111111111111110111","111111111111110100","111111111111110100","000000000000001001","111111111111101011","111111111111111110","000000000000010010","111111111111111111","111111111111111001","000000000000000010","111111111111101110","000000000000011000","000000000000000000","000000000000000000","000000000000110100","000000000000010101","111111111111001111","111111111111011101","000000000000000010","111111111111111111","000000000000010110","000000000000000101"),
("000000000000000110","000000000000001001","111111111111110001","111111111111100010","111111111111110100","000000000000011100","111111111111010101","000000000000101000","111111111111001101","111111111111101101","000000000000011010","000000000000001011","111111111111111101","000000000000001100","111111111111100110","000000000000000001","000000000000011101","111111111111111010","111111111111111011","111111111111111011","111111111111100010","000000000000000101","000000000000000011","000000000000000000","000000000000001101","111111111111100111","000000000000011100","111111111111101010","111111111111010011","111111111111111000","111111111111111101","111111111111100110","111111111111100001","111111111111111100","000000000000000010","000000000000000010","111111111111111010","111111111111110011","000000000000000010","000000000000000110","111111111111101001","000000000000010001","000000000000001100","111111111111110110","000000000000001110","111111111111111110","000000000000000011","000000000000000011","000000000000011100","000000000000001001","000000000000010001","000000000000101001","111111111111100101","111111111111111010","111111111111110001","000000000000010010","000000000000011000","111111111111100110","111111111111111111","000000000000000001","111111111111111001","111111111111111011","111111111111000111","000000000000010101","111111111111000101","000000000000010000","111111111111111010","000000000000010000","000000000000001011","000000000000000010","000000000000001000","111111111111111101","111111111111111000","111111111111011000","111111111111111110","111111111111111110","111111111111110111","111111111111110110","000000000000001001","000000000000100000","000000000000010000","000000000000000001","111111111111111000","111111111111111111","111111111111111001","000000000000000110","111111111111111111","000000000000000000","000000000000000011","111111111111110110","000000000000011001","000000000000010101","111111111110100110","111111111111010111","111111111111110011","111111111111110101","111111111111011110","111111111111010011","111111111111110011","000000000000001111","111111111111111110","000000000000100100","111111111111111101","000000000000100101","111111111111110000","000000000000001010","111111111111110010","111111111111111101","111111111111110111","000000000000000001","111111111111110011","111111111111101010","000000000000001010","000000000000010001","000000000000101101","111111111111111101","111111111111101111","111111111111110111","000000000000001010","000000000000000000","000000000000101010","111111111111101110","111111111111010111","111111111111110110","111111111111111101","111111111111111100","111111111111111011","000000000000000010"),
("000000000000100100","111111111111101000","000000000000001100","111111111111001010","000000000000000101","000000000000000100","111111111111100101","111111111111101100","111111111111010101","111111111111110001","111111111111110011","000000000000101111","000000000000000000","111111111111101110","111111111111110001","111111111111110101","000000000000000010","111111111111110010","000000000000001010","111111111111011100","111111111111011110","111111111111111011","111111111111011011","000000000000000000","000000000000001000","111111111111110010","000000000000000110","111111111111010001","111111111111101001","000000000000100001","000000000000000101","111111111111101110","111111111111100111","000000000000101010","000000000000010000","111111111111110011","000000000000000101","000000000000001110","000000000000000011","000000000000001011","000000000000010011","000000000000110110","000000000000001010","111111111111011010","000000000000100110","111111111111110100","111111111111111001","111111111111111111","000000000000010101","000000000000000101","111111111111011100","000000000000011000","111111111111101100","000000000000000111","000000000000000010","111111111111101110","000000000000100100","111111111111100011","111111111111110110","111111111111111001","111111111111111011","111111111111101100","111111111110010011","111111111111110000","111111111111111000","111111111111111100","000000000000010100","000000000000100101","000000000000011011","111111111111111000","111111111111111010","111111111111111011","000000000000010100","111111111111011111","000000000000001000","111111111111101101","000000000000000000","111111111111011110","111111111111101001","111111111111110110","000000000000000111","000000000000011010","111111111111101101","111111111111100110","111111111111110110","111111111111110100","000000000000010000","000000000000100001","111111111111110010","111111111111111101","000000000000101000","111111111111111101","111111111111010110","111111111111001001","111111111111110000","111111111111100011","111111111111011010","000000000000000101","000000000000011101","000000000000010100","000000000000000000","000000000000010011","000000000000010000","000000000000001111","000000000000000000","000000000000000000","111111111111110000","111111111111111000","111111111111111010","111111111111011101","000000000000000000","111111111111111100","000000000000111101","000000000000010101","000000000000010100","111111111111101111","000000000000000000","000000000000011110","111111111111110110","111111111111111001","000000000000100111","000000000000001011","111111111111010001","111111111111111101","111111111111101000","111111111111111011","000000000000100011","000000000000011001"),
("000000000001000100","111111111111100001","000000000000010011","111111111111101000","000000000000001000","000000000000000001","111111111111100010","111111111111110101","000000000000000101","111111111111000110","111111111111011110","000000000000111000","000000000000000110","111111111111011011","111111111111011000","111111111111101111","111111111111110111","000000000000000011","000000000000010101","111111111111101101","111111111111101110","111111111111101101","111111111111101001","111111111111111100","000000000000011111","000000000000000100","000000000000001001","111111111111110101","000000000000010001","000000000000001111","000000000000101111","111111111111111000","111111111111110100","000000000000100101","000000000000101111","000000000000001000","000000000000010011","000000000000011101","111111111111110001","000000000000001100","000000000000101111","000000000000101111","000000000000001000","111111111111100011","000000000000101100","111111111111110111","000000000000000011","000000000000100110","000000000000011000","000000000000100010","111111111111011010","000000000000001010","111111111111100101","000000000000100111","000000000000000011","111111111111101100","000000000000110110","111111111111001101","111111111111010101","111111111111111010","000000000000010100","111111111111101010","111111111110101101","111111111111101111","111111111111000110","000000000000000110","000000000000011111","000000000000001111","111111111111111011","111111111111111001","000000000000001100","000000000000001111","000000000000000011","111111111111101110","000000000000000000","111111111111110111","000000000000100101","111111111111100101","111111111111101001","000000000000000000","111111111111110101","000000000000100000","111111111111101001","111111111111011000","111111111111110010","111111111111101100","000000000001000001","000000000000101000","111111111111101110","111111111111110101","000000000000010010","000000000000000000","111111111111101100","111111111110111110","111111111111100000","000000000000001010","111111111111111111","000000000000011010","000000000000010111","000000000000000110","000000000000110101","000000000000011100","111111111111101110","000000000000000111","111111111111110110","111111111111110000","111111111111110010","111111111111011100","111111111111110000","111111111111100100","000000000000010011","111111111111110110","000000000000011111","000000000000000000","000000000000000000","111111111111101011","000000000000000001","000000000000101000","111111111111101010","000000000000101100","000000000001011011","000000000000000111","000000000000001100","111111111111010000","111111111111101100","111111111111111101","000000000000111011","111111111111110101"),
("000000000000011000","000000000000010001","000000000000100000","111111111111111011","000000000000010010","111111111111111111","111111111111110100","111111111111110100","111111111111110111","111111111111100011","111111111111101110","000000000000001111","111111111111110011","111111111111111110","111111111111110011","000000000000000011","111111111111111010","000000000000000101","000000000000001011","111111111111110011","000000000000000000","000000000000000001","111111111111011001","111111111111100000","000000000000000001","000000000000000000","000000000000010100","111111111111100100","000000000000000000","000000000000011001","000000000000000101","000000000000000000","000000000000000011","000000000000100001","000000000000001001","000000000000000000","000000000000011000","000000000000000101","000000000000001000","000000000000100100","000000000000001011","000000000000011000","111111111111111101","000000000000001011","000000000000011110","111111111111111110","111111111111111001","111111111111111101","000000000000100110","000000000000001000","111111111111001100","111111111111110111","111111111111101110","000000000000001011","111111111111110110","111111111111111101","000000000000011011","111111111111110011","111111111111011001","000000000000001111","000000000000001110","111111111111111011","111111111111101111","111111111111111101","111111111111101010","000000000000001010","000000000000000110","000000000000010011","111111111111111001","000000000000011101","000000000000000100","111111111111111001","000000000000000011","000000000000000000","111111111111110111","111111111111111010","000000000000100011","111111111111011100","111111111111101101","000000000000000001","000000000000100000","000000000000011100","111111111111110001","000000000000001101","111111111111111111","111111111111110000","000000000000011001","000000000000101110","111111111111110111","111111111111110110","111111111111111010","111111111111110001","000000000000000000","111111111111001101","111111111111110101","111111111111110101","000000000000000000","111111111111110110","000000000000001001","000000000000010011","000000000000101001","000000000000010000","111111111111111110","111111111111100110","111111111111111101","000000000000000010","000000000000000000","111111111111111010","111111111111110101","111111111111101000","111111111111111000","111111111111111011","000000000000001001","000000000000000101","000000000000000011","111111111111110111","000000000000001010","000000000000001111","000000000000010101","000000000000100101","000000000000100100","000000000000000011","111111111111110111","111111111111011100","000000000000000001","000000000000000100","000000000000000011","000000000000100010"),
("000000000000000100","000000000000001001","000000000000010110","111111111111101111","000000000000000000","000000000000000010","000000000000010000","111111111111101101","111111111111100100","111111111111011001","111111111111111010","000000000000010011","000000000000000111","111111111111011111","000000000000000010","111111111111111011","000000000000000001","111111111111101011","111111111111101001","111111111111101101","111111111111110011","111111111111111111","111111111111110001","111111111111010100","111111111111110000","000000000000101000","111111111111100010","000000000000000111","000000000000010010","000000000000001001","000000000000001000","111111111111101011","111111111111100000","000000000000010111","000000000000001000","000000000000000000","111111111111111101","111111111111110010","111111111111100100","000000000000001011","111111111111110100","000000000000001100","111111111111111101","000000000000001000","111111111111111011","111111111111111101","000000000000001101","000000000000000111","000000000000000110","000000000000000010","111111111111101110","111111111111100000","000000000000000000","000000000000100100","111111111111101010","000000000000000001","111111111111111111","111111111111110110","111111111111100101","111111111111110100","111111111111100111","111111111111011101","111111111111111100","000000000000001110","111111111111111000","111111111111100011","111111111111101101","000000000000100101","000000000000000100","111111111111101111","000000000000001001","111111111111110000","000000000000001111","111111111111110001","111111111111101101","111111111111101111","000000000000001101","000000000000001111","000000000000010101","000000000000001011","111111111111111101","000000000000000111","000000000000010100","000000000000011100","111111111111101100","111111111111010000","000000000000000000","111111111111110100","000000000000001111","111111111111111011","111111111111101011","000000000000000100","000000000000010100","111111111111111010","111111111111111010","111111111111110010","000000000000001110","000000000000000010","111111111111111100","000000000000001010","000000000000011111","000000000000001111","000000000000010100","111111111111100111","111111111111111101","111111111111111100","111111111111101010","111111111111111110","111111111111110111","000000000000000000","111111111111101000","111111111111110101","000000000000011011","000000000000000001","111111111111111101","000000000000010101","000000000000010010","000000000000100000","111111111111110000","000000000000110001","000000000000001000","111111111111111110","000000000000010001","000000000000010000","000000000000000000","000000000000000111","111111111111111110","111111111111110010"),
("000000000000001101","111111111111110101","000000000000000100","111111111111111100","111111111111110101","000000000000000000","000000000000010010","111111111111110011","000000000000010001","111111111111110110","000000000000001101","111111111111101100","111111111111111101","000000000000010100","000000000000001101","000000000000001110","000000000000000111","111111111111110100","000000000000000101","111111111111110111","000000000000000100","111111111111110001","000000000000001000","111111111111101110","000000000000001110","111111111111110110","000000000000010000","111111111111101101","111111111111110011","000000000000000110","111111111111110000","111111111111101101","111111111111111001","000000000000010010","111111111111110011","111111111111110110","000000000000001011","000000000000001111","111111111111110010","111111111111101101","000000000000001011","111111111111101111","000000000000000000","111111111111111001","111111111111101111","111111111111101101","111111111111111101","111111111111111111","000000000000000001","111111111111101110","000000000000000000","000000000000000000","111111111111111111","111111111111111110","111111111111110001","000000000000001101","111111111111110011","111111111111101111","000000000000000100","000000000000010010","000000000000000100","111111111111111010","000000000000001101","000000000000001000","111111111111111001","000000000000001111","000000000000001000","111111111111111101","111111111111111110","000000000000000000","000000000000000100","111111111111101101","000000000000001001","111111111111111111","111111111111110000","111111111111110010","000000000000010000","000000000000000001","000000000000001000","111111111111110101","000000000000001010","000000000000001101","000000000000010010","111111111111111001","111111111111111110","111111111111101101","111111111111111010","000000000000010000","000000000000001110","000000000000000001","000000000000000001","000000000000001100","000000000000000111","111111111111110000","111111111111111101","000000000000001010","111111111111111001","111111111111111101","000000000000001010","000000000000001001","000000000000010001","000000000000001111","000000000000000000","000000000000010011","111111111111110011","000000000000001101","111111111111110110","111111111111111100","000000000000000100","000000000000010100","000000000000000010","111111111111101110","111111111111111101","000000000000001100","111111111111111000","000000000000001000","111111111111111111","111111111111111000","111111111111111000","111111111111101100","111111111111110101","111111111111110110","000000000000001111","111111111111110000","000000000000010010","111111111111110101","111111111111110000","000000000000001001"),
("111111111111011100","111111111111110101","111111111111101010","000000000000001101","000000000000001111","111111111111111010","111111111111110000","111111111111100111","000000000000100001","000000000000101110","000000000000010100","000000000000010000","000000000000010110","111111111111110010","111111111111111111","000000000000010011","000000000000100000","000000000000010100","000000000000001110","000000000000010100","111111111111101100","000000000000010101","000000000000001110","111111111111100011","111111111111110110","111111111111111010","000000000000000000","000000000000000010","000000000000011001","000000000000001001","111111111111100101","000000000000100011","000000000000011011","111111111111001111","111111111111111101","111111111111110101","111111111111101111","000000000000000000","111111111111110110","000000000000100001","000000000000000110","111111111111100110","000000000000011110","111111111111101110","111111111111100101","000000000000100100","000000000000010010","111111111111110011","000000000000011101","000000000000011110","000000000000011001","111111111111111100","000000000000000011","111111111111111001","000000000000011010","000000000000000111","111111111111110111","000000000000010000","000000000000000101","000000000000001000","000000000000100110","000000000000100100","000000000000100111","111111111111100111","111111111111100001","111111111111111011","111111111111010011","000000000000001011","000000000000011010","000000000000001001","000000000000010110","000000000000100001","111111111111111001","000000000000100110","000000000000001110","000000000000000110","111111111111100011","000000000000100100","111111111111110111","000000000000001110","111111111111011001","111111111111110100","111111111111101100","000000000000100011","000000000000011110","111111111111111000","000000000000001101","000000000000000000","111111111111110001","000000000000000010","111111111111101001","111111111111111111","000000000000000100","111111111111111111","000000000000000000","111111111111100111","000000000000010000","000000000000010000","000000000000001111","000000000000110100","111111111111111100","000000000000000101","000000000000000111","111111111111111000","000000000000000110","000000000000000100","111111111111110101","000000000000000101","000000000000000010","111111111111100101","111111111111110101","111111111111011100","000000000000000110","000000000000100100","000000000000010111","111111111111111011","000000000000011000","000000000000100101","111111111111011000","000000000000000001","000000000000001111","111111111111111101","111111111111111001","000000000000001100","000000000000000110","111111111111100001","111111111111111010","000000000000000010"),
("000000000000000001","111111111111011111","000000000000001100","111111111111111010","111111111111011011","111111111111011110","111111111111111100","111111111111110001","000000000000010100","000000000000000001","111111111111100010","000000000000000100","000000000000010110","000000000000001101","000000000000011010","000000000000010001","111111111111110100","000000000000000010","000000000000010101","000000000000101101","000000000000001000","000000000000100111","111111111111100111","000000000000001011","000000000000010100","111111111111110000","111111111111011101","000000000000000101","000000000000000001","000000000000000100","000000000000001001","111111111111111101","111111111111110000","111111111111101100","000000000000001000","111111111111101110","000000000000101111","111111111111111011","111111111111101110","000000000000001010","111111111111110101","111111111111100101","000000000000101000","111111111111011001","111111111111100101","111111111111110101","000000000000000111","111111111111110000","000000000000001110","000000000000000101","000000000000000101","111111111111100110","111111111111111100","000000000000000100","000000000000110111","000000000000100101","111111111111101001","000000000000001011","000000000000010000","111111111111110111","000000000000000011","000000000000100101","111111111111110101","000000000000000000","111111111111100000","000000000000110010","111111111111110111","111111111111111100","000000000000011010","000000000000010011","111111111111100111","111111111111111001","111111111111101101","000000000000001110","111111111111111101","000000000000001101","111111111111110100","000000000000010010","000000000000010100","000000000000101011","111111111111010000","111111111111100010","111111111111101001","000000000000011100","111111111111101010","000000000000010010","000000000000101110","111111111111110100","111111111111111011","000000000000001110","000000000000000111","111111111111110010","000000000000111011","111111111111111011","000000000000010101","000000000000000000","000000000000001111","000000000000001001","111111111111110111","000000000000010110","111111111111111110","111111111111101011","111111111111101111","111111111111100011","111111111111110101","111111111111011110","000000000000010000","000000000000100111","000000000000001010","000000000000101101","111111111111111011","111111111111110111","111111111111100101","000000000000010011","000000000000101001","111111111111110111","111111111111111011","000000000000010100","000000000000010011","000000000000000011","000000000000011001","000000000000001011","111111111111101110","000000000000110010","000000000000000000","111111111111101010","000000000000100001","111111111111110011"),
("111111111111110101","111111111111100011","000000000000011000","111111111111110011","000000000000010101","111111111111110011","000000000000001000","000000000000000000","000000000000100000","000000000000001101","000000000000010011","111111111111010010","000000000000001000","000000000000001101","000000000000100000","000000000000000000","000000000000100110","111111111111111001","000000000000100010","000000000000011111","000000000000010001","000000000000010101","000000000000011001","111111111111110011","000000000000010010","111111111111100110","000000000000000000","000000000000000111","000000000000111101","111111111111110111","111111111111100101","000000000000000000","000000000000010100","111111111111010110","111111111111110101","000000000000000010","111111111111111101","111111111111111110","111111111111110000","000000000000100000","000000000000000111","111111111111010100","000000000000010001","000000000000000101","111111111111111000","000000000000010110","000000000000001101","111111111111101000","000000000000000010","111111111111101010","000000000000001011","000000000000000000","111111111111101100","000000000000001111","000000000000101001","000000000000010110","111111111111100011","000000000000010000","000000000000011000","000000000000001110","111111111111111000","000000000000000101","000000000000000011","000000000000000000","111111111111110101","111111111111111110","000000000000000001","111111111111111101","000000000000000110","000000000000000101","000000000000000101","000000000000001011","000000000000011101","000000000000111001","111111111111100110","000000000000001110","000000000000000000","000000000000000010","000000000000001100","000000000000101001","111111111111100001","111111111111100100","000000000000001110","000000000000101010","000000000000000011","000000000000001011","000000000000100011","000000000000000101","111111111111100101","111111111111111111","111111111111011110","111111111111100100","111111111111110110","111111111111111000","000000000000010000","000000000000001110","111111111111111001","000000000000010110","111111111111110001","000000000000010010","000000000000000000","111111111111011010","111111111111100111","111111111111100101","000000000000001111","111111111111101100","000000000000000001","000000000000000000","111111111111100101","000000000000001000","000000000000010000","111111111111101010","111111111111111110","000000000000000100","000000000000001000","111111111111111011","000000000000000101","000000000000000111","111111111111100110","000000000000100010","000000000000010000","111111111111101100","111111111111100011","000000000000110101","111111111111110110","111111111111010001","000000000000001000","000000000000000000"),
("111111111111011111","111111111111101110","111111111111110011","000000000000001100","000000000000011100","000000000000001000","111111111111101110","000000000000001100","000000000000110001","000000000000101100","000000000000000111","000000000000000000","000000000000010110","111111111111110011","000000000000010101","000000000000010011","000000000000110111","000000000000000100","000000000000011100","000000000000001001","000000000000000000","000000000000110001","111111111111111111","000000000000000000","000000000000000110","000000000000000100","111111111111110100","111111111111111111","000000000000101010","000000000000000101","111111111111000110","000000000000000000","111111111111111000","111111111111000011","111111111111010011","000000000000000010","111111111111100011","000000000000000010","111111111111111101","111111111111111110","111111111111100110","111111111111011000","000000000000100110","000000000000010100","000000000000010111","111111111111111110","000000000000111001","111111111110111000","000000000000000101","111111111111110000","000000000000101010","000000000000010111","111111111111110011","111111111111100011","000000000000000010","000000000000000111","111111111111010100","000000000000010011","111111111111011011","000000000000010001","111111111111101000","000000000000000100","000000000000000010","111111111111101110","111111111111111011","111111111111100111","000000000000011010","000000000000010001","000000000000100110","000000000000001101","000000000000000000","000000000000000101","000000000000100011","000000000000100010","000000000000011101","000000000000001000","111111111111100100","000000000000001111","111111111111111111","000000000000101101","111111111111101100","111111111111011000","000000000000100100","111111111111110000","000000000000000010","000000000000011000","000000000000000010","000000000000100100","000000000000000011","000000000000001000","111111111111110100","111111111111100101","111111111111110110","000000000000000010","111111111111101000","111111111111101010","000000000000001010","000000000000010100","111111111111111010","111111111111100101","111111111111100100","111111111111100000","111111111111100111","000000000000001100","000000000000010011","000000000000001110","111111111111110101","000000000000010101","000000000000010000","111111111111111101","111111111111111110","000000000000010000","000000000000101001","000000000000100111","111111111111011010","000000000000001111","000000000000000011","000000000000001110","111111111111001111","000000000000010001","111111111111110010","111111111111111010","111111111111100010","000000000000100110","000000000000000001","111111111111001101","000000000000000000","111111111111110100"),
("111111111111011000","111111111111111100","111111111111110100","111111111111101111","000000000001000110","111111111111101110","111111111111100001","000000000000011001","000000000000010011","000000000000010110","111111111111111100","000000000000001101","111111111111100010","111111111111100111","000000000000001011","000000000000001001","000000000000101000","000000000000010011","000000000000100010","000000000000010000","111111111111101000","111111111111111011","000000000000010001","111111111111110101","111111111111101101","111111111111101011","000000000000111000","111111111111101100","000000000000101111","111111111111011111","111111111111010111","111111111111110111","000000000000010011","111111111111100111","111111111111110010","000000000000001110","000000000000010000","000000000000100101","111111111111111100","000000000000010101","111111111111111010","111111111111010101","000000000000001000","111111111111111000","000000000000000000","000000000000001000","000000000000011111","111111111111100110","000000000000100101","111111111111110110","000000000000010010","000000000000101011","111111111111101101","111111111111001011","000000000000001000","111111111111110100","111111111111010011","111111111111111010","111111111111101100","111111111111111101","111111111111111000","111111111111111100","000000000000010101","111111111111111111","111111111111100100","111111111111110100","000000000000000011","111111111111110001","000000000000001100","111111111111110000","111111111111100010","000000000000000101","000000000000001000","111111111111110111","111111111111111110","000000000000100000","111111111111111110","111111111111111010","111111111111111010","000000000000001010","111111111111110101","111111111111100100","111111111111111010","111111111111000110","000000000000010001","000000000000001011","000000000000101100","000000000000110110","111111111111100110","111111111111110110","111111111111111100","111111111111101111","000000000000000000","111111111111111100","111111111111110101","111111111111001111","000000000000001001","000000000000001001","111111111111011011","111111111111110010","111111111111100100","111111111111100111","111111111111011011","111111111111111000","111111111111101100","000000000000001111","111111111111101010","111111111111110111","111111111111101100","000000000000011000","111111111111101100","000000000000000000","000000000000001001","000000000000000101","000000000000001000","111111111111101000","000000000000010100","000000000000001010","111111111111011010","000000000000000100","111111111111100111","111111111111011010","111111111111110100","000000000000001100","000000000000011111","111111111111010011","000000000000001110","111111111111110100"),
("111111111110110100","000000000000000010","111111111111111011","111111111111100111","000000000000011100","111111111111101100","000000000000000000","000000000000011001","000000000000010010","111111111111111101","111111111111110011","000000000000010000","000000000000001001","111111111111101110","000000000000001011","000000000000000101","000000000000010001","000000000000010011","000000000000110001","000000000000001110","000000000000000101","111111111111101111","000000000000000011","000000000000011000","111111111111111111","111111111111101101","000000000000011010","000000000000001010","000000000000101011","111111111111100111","111111111111011001","111111111111101100","000000000000000111","111111111111011010","000000000000000011","000000000000010101","000000000000100011","000000000000001100","111111111111110111","000000000000000000","000000000000010101","111111111111010011","000000000000000111","111111111111111111","111111111111110111","000000000000000000","000000000000000111","111111111111100001","000000000000101100","000000000000010010","000000000000011111","000000000000011011","000000000000000000","000000000000001111","000000000000010010","111111111111111110","111111111111101100","000000000000001011","000000000000011101","000000000000000000","111111111111110110","000000000000001101","000000000000010011","111111111111010111","111111111111001101","000000000000000101","111111111111100011","111111111111011011","000000000000001000","000000000000010011","111111111111011111","111111111111111001","111111111111111111","000000000000001010","111111111111110010","000000000000010010","111111111111100111","111111111111110111","000000000000001110","000000000000000001","111111111111101110","111111111111011101","111111111111100100","111111111111010001","111111111111111111","000000000000011101","000000000000100100","111111111111111010","111111111111010110","000000000000011111","111111111111010111","111111111111111010","111111111111110000","111111111111110000","111111111111110011","111111111111101101","000000000000001011","000000000000001111","111111111111101000","111111111111101101","111111111111100010","111111111111101110","111111111111011000","111111111111110001","111111111111100110","111111111111110001","000000000000001001","000000000000100101","111111111111111101","000000000000000101","000000000000011001","000000000000000110","111111111111100010","000000000000000010","111111111111110101","111111111111100010","111111111111111011","111111111111111111","111111111111011010","000000000000011100","000000000000001011","111111111111100001","000000000000000000","000000000000000101","000000000000000101","111111111111011000","000000000000101000","111111111111111100"),
("111111111111011011","000000000000001001","111111111111111110","111111111111111000","000000000000100000","111111111111101010","111111111111110010","000000000000010011","000000000000011010","000000000000000010","000000000000000000","000000000000110010","000000000000000101","111111111111100000","000000000000011110","000000000000000011","111111111111111010","000000000000011101","000000000000000100","000000000000010010","111111111111101100","000000000000000010","111111111111101110","000000000000000100","111111111111100011","111111111111110011","000000000000001010","111111111111101000","000000000000000001","111111111111011110","111111111111100010","111111111111110100","111111111111110101","111111111111100001","111111111111111001","111111111111111100","000000000000010001","000000000000001101","111111111111101001","000000000000010111","000000000000000011","111111111111011100","000000000000001011","000000000000010001","111111111111111000","000000000000010010","000000000000001100","111111111111110000","000000000000011011","111111111111110011","000000000000001011","111111111111110010","000000000000010000","000000000000010000","000000000000000100","111111111111111110","111111111111010110","000000000000010001","000000000000001010","111111111111111010","111111111111111011","000000000000010111","000000000000010001","111111111111101110","111111111111000010","000000000000001111","000000000000000000","111111111111101011","000000000000001001","000000000000001101","111111111111100011","111111111111111101","111111111111110001","000000000000001000","000000000000001011","111111111111101111","000000000000001101","000000000000001001","000000000000010000","000000000000001100","111111111111100000","111111111111110000","111111111111001110","000000000000000110","000000000000001100","111111111111100101","000000000000100010","111111111111110101","111111111111101101","111111111111111100","111111111111001110","111111111111101100","000000000000100011","111111111111111011","111111111111111100","111111111111011111","111111111111110111","000000000000010101","111111111111100010","111111111111110010","111111111111000110","000000000000010001","111111111111101010","111111111111111110","111111111111111011","111111111111111010","111111111111101111","000000000000010011","000000000000010111","111111111111110001","111111111111111011","111111111111110101","111111111111111110","000000000000010101","000000000000010001","111111111111011000","111111111111111100","000000000000001001","111111111111010000","000000000000101011","000000000000010010","111111111111101110","111111111111110110","000000000000000100","000000000000000000","111111111111011000","000000000000000110","000000000000000110"),
("111111111111010101","111111111111110011","111111111111111111","000000000000000011","000000000000010000","111111111111011110","000000000000000000","000000000000110111","000000000000000011","111111111111101000","000000000000000111","000000000000010001","000000000000011001","111111111111111110","000000000000010000","000000000000011011","111111111111100100","111111111111111101","111111111111101111","000000000000001110","111111111111100100","111111111111110111","111111111111011110","111111111111001110","111111111111111110","000000000000001000","000000000000010000","000000000000011001","111111111111101011","111111111111100110","111111111111111010","111111111111101111","000000000000000010","111111111111011100","111111111111111100","000000000000011000","000000000000010111","111111111111110101","000000000000000100","000000000000010000","000000000000010101","111111111111110110","000000000000001000","111111111111110101","000000000000001101","111111111111101010","111111111111100010","000000000000000100","000000000000011010","000000000000000110","111111111111110101","000000000000001011","111111111111110100","000000000000101111","000000000000000111","111111111111111100","111111111111111011","000000000000010101","111111111111110100","111111111111110011","111111111111111101","000000000000010001","111111111111111001","111111111111111110","111111111111101011","111111111111110111","111111111111100100","111111111111101011","000000000000001000","111111111111100100","111111111111110111","000000000000000000","111111111111011101","111111111111100101","000000000000001110","000000000000001011","000000000000011000","000000000000010001","000000000000001011","000000000000001011","111111111111101010","000000000000000010","111111111111100000","111111111111111011","000000000000001101","111111111111101101","000000000000001101","000000000000001010","111111111111111111","111111111111101001","111111111111110100","111111111111110101","000000000000100100","111111111111001101","000000000000000000","111111111111001101","000000000000100011","000000000000110100","111111111111100101","111111111111111111","111111111111101000","000000000000100010","111111111111101101","000000000000001011","111111111111101101","111111111111110000","000000000000001111","000000000000001101","111111111111110111","111111111111110010","000000000000000101","000000000000000101","000000000000000100","000000000000000010","000000000000000010","111111111111011110","000000000000010101","111111111111110111","111111111111100101","000000000000101101","000000000000010100","111111111111101000","000000000000010100","000000000000011001","111111111111101010","111111111111101101","000000000000001010","111111111111111110"),
("111111111111000011","111111111111111001","111111111111111101","111111111111111001","000000000000011111","111111111111011110","000000000000000000","000000000000100111","000000000000001101","000000000000000101","111111111111100100","000000000000011001","000000000000011001","000000000000001100","000000000000001101","000000000000011000","111111111111111011","000000000000001011","000000000000010011","000000000000000001","111111111111011100","111111111111011110","111111111111110101","111111111111100010","000000000000000000","111111111111100111","000000000000001101","000000000000000000","111111111111110111","111111111111111010","111111111111101000","111111111111111001","000000000000001101","000000000000000000","000000000000000010","111111111111110110","000000000000010001","111111111111100111","000000000000000000","111111111111110001","000000000000000111","000000000000010000","111111111111111110","111111111111110000","111111111111110011","111111111111101110","111111111111110011","000000000000010111","000000000000010111","000000000000011101","000000000000010111","000000000000000101","000000000000000001","000000000000100110","000000000000010100","000000000000001011","000000000000000111","111111111111110101","000000000000000000","000000000000000010","111111111111100100","000000000000010110","000000000000010000","111111111111101111","111111111111100110","000000000000011001","111111111111010110","111111111111101001","000000000000001111","000000000000010011","111111111111101101","000000000000011001","111111111111100000","111111111111111101","111111111111111011","000000000000001010","000000000000000000","000000000000000001","111111111111111010","000000000000011000","111111111111011111","111111111111111011","111111111111110010","000000000000101010","000000000000000010","000000000000000111","111111111111111100","000000000000000001","111111111111111111","000000000000010000","111111111111111110","111111111111110010","000000000000010011","111111111111111011","000000000000100000","111111111111001001","000000000000011101","000000000000010000","111111111111101010","111111111111100011","111111111111011111","000000000000011110","111111111111101101","000000000000000000","111111111111100011","111111111111111011","000000000000000101","111111111111111101","000000000000000110","000000000000001011","111111111111110100","000000000000010100","000000000000010001","111111111111111011","000000000000000010","111111111111100101","111111111111111100","000000000000000010","111111111111110010","000000000000000111","000000000000001000","000000000000000011","000000000000001110","111111111111111111","000000000000000110","000000000000010010","000000000000100110","000000000000010011"),
("111111111111001000","000000000000010011","000000000000001100","111111111111110001","111111111111011100","111111111111110101","000000000000000011","000000000000001101","000000000000000011","000000000000001011","111111111111101011","000000000000101100","000000000000101000","111111111111100010","000000000000001010","000000000000010110","111111111111111110","000000000000001101","111111111111111000","000000000000011000","111111111111111011","111111111111111111","111111111111110011","111111111111111100","000000000000001011","000000000000001011","000000000000011101","000000000000010011","000000000000001110","111111111111110011","000000000000001011","000000000000001001","000000000000001110","000000000000000111","000000000000001010","111111111111111100","000000000000001101","111111111111110100","000000000000011110","000000000000000000","000000000000001000","000000000000000101","000000000000001110","111111111111101011","000000000000010001","111111111111111010","111111111111101110","000000000000000001","000000000000000111","111111111111110001","000000000000011101","000000000000000110","000000000000001110","000000000000100101","000000000000010011","111111111111111001","000000000000011110","111111111111111001","000000000000010101","000000000000001011","000000000000000010","000000000000010110","000000000000011100","111111111111101101","111111111111010001","000000000000100010","111111111111001001","111111111111101000","000000000000010100","000000000000001101","000000000000001000","000000000000001110","111111111111100001","000000000000001111","111111111111111100","111111111111110011","111111111111110110","000000000000000001","111111111111111111","000000000000010001","000000000000000000","000000000000001100","000000000000000000","000000000000111011","111111111111110110","111111111111101011","000000000000001001","000000000000000110","000000000000000000","111111111111110001","000000000000100000","111111111111111000","000000000000011100","111111111111110100","111111111111111011","111111111111110111","000000000000001110","000000000000001010","111111111111100011","111111111111100110","111111111111011101","000000000000100110","111111111111001001","111111111111101111","000000000000010010","111111111111110001","000000000000000010","000000000000010110","000000000000001101","111111111111110111","111111111111111011","000000000000000001","000000000000001011","111111111111110011","111111111111111000","111111111111011111","000000000000000001","000000000000010110","000000000000001001","000000000000001110","000000000000010011","000000000000010110","111111111111110010","111111111111111011","000000000000001110","000000000000101000","000000000000010001","000000000000001110"),
("111111111111111001","000000000000011100","111111111111110011","111111111111111010","111111111110101110","111111111111101001","000000000000010011","111111111111111100","111111111111110110","000000000000010110","000000000000000011","000000000000000101","000000000000010110","111111111111111100","111111111111111101","000000000000010001","000000000000001011","000000000000000111","111111111111110110","000000000000010010","111111111111101110","111111111111111010","000000000000000010","000000000000000000","000000000000000110","111111111111110001","000000000000000001","000000000000001110","000000000000000001","000000000000000110","111111111111111011","111111111111101011","000000000000001100","111111111111111010","111111111111101111","111111111111101101","000000000000000100","111111111111101111","000000000000100010","111111111111110010","000000000000001001","000000000000010101","000000000000010001","000000000000001011","111111111111111001","111111111111110110","111111111111100001","000000000000000000","000000000000000000","000000000000010001","000000000000001100","000000000000000001","111111111111111101","000000000000011010","000000000000010010","111111111111111010","000000000000001110","111111111111111010","000000000000001011","111111111111111010","111111111111010010","000000000000010000","000000000000001000","000000000000000011","111111111111110011","000000000000000000","111111111111001111","000000000000000101","000000000000010101","000000000000011100","111111111111101011","000000000000010000","111111111111100101","111111111111101011","111111111111111001","000000000000000110","000000000000010000","000000000000010100","000000000000000000","000000000000010110","111111111111110010","000000000000010100","111111111111101110","000000000000100100","111111111111111001","000000000000001100","111111111111111101","000000000000000110","000000000000001011","111111111111111111","000000000000010011","000000000000000101","111111111111111010","111111111111110111","111111111111110111","111111111111111011","000000000000001010","000000000000001111","111111111111110110","000000000000001100","111111111111111111","111111111111111101","111111111111010111","000000000000000110","000000000000010111","000000000000001110","000000000000000100","000000000000000101","111111111111111011","111111111111111000","111111111111111101","000000000000011101","000000000000000010","111111111111111001","000000000000000100","111111111111100111","000000000000000111","000000000000010010","000000000000100011","000000000000011000","000000000000100001","000000000000010101","000000000000001101","111111111111111001","000000000000000000","000000000000101011","000000000000001101","000000000000010111"),
("111111111111011110","000000000000100000","111111111111111100","000000000000001100","111111111110100110","111111111111111000","000000000000000110","000000000000001111","111111111111111000","111111111111111011","111111111111100111","000000000000001010","000000000000100101","111111111111110111","000000000000001110","000000000000100010","111111111111101101","000000000000001001","000000000000000101","000000000000010010","111111111111111110","111111111111111100","000000000000010010","000000000000010100","000000000000001111","000000000000010000","111111111111110111","000000000000100110","000000000000000000","000000000000001010","000000000000000100","000000000000000011","111111111111110101","000000000000010111","000000000000000101","111111111111111010","000000000000011010","111111111111110011","000000000000001111","000000000000001000","111111111111111011","000000000000001101","000000000000001000","111111111111110000","111111111111111000","111111111111110100","000000000000000000","111111111111110101","111111111111110101","000000000000000010","000000000000010010","111111111111100101","000000000000001100","000000000000110011","000000000000001100","000000000000000001","000000000000011000","000000000000001110","000000000000011010","111111111111110011","111111111111101110","111111111111111111","000000000000010100","111111111111100110","111111111111111110","111111111111111100","111111111111101001","111111111111111111","000000000000010010","000000000000010111","000000000000001001","000000000000100001","111111111111001010","111111111111111010","000000000000010010","000000000000001001","000000000000000010","000000000000001110","111111111111110000","000000000000000111","111111111111111111","000000000000010100","111111111111101001","000000000000000000","000000000000011001","111111111111110010","111111111111101001","111111111111011110","111111111111111010","111111111111111011","000000000000001100","000000000000000001","111111111111111001","111111111111101100","000000000000011101","111111111111110100","111111111111100111","000000000000001011","111111111111111111","000000000000010001","111111111111100101","111111111111110101","111111111111110011","111111111111110000","000000000000010010","111111111111110100","000000000000000000","111111111111111001","000000000000001110","000000000000000010","000000000000010100","000000000000011110","000000000000000011","000000000000000011","111111111111111111","111111111111011000","111111111111111111","000000000000000111","000000000000000100","000000000000101011","000000000000101101","000000000000001111","000000000000011011","000000000000000010","111111111111110101","000000000000011110","000000000000000111","000000000000001101"),
("111111111111111110","000000000000011111","000000000000010001","000000000000001111","111111111110011101","000000000000000000","000000000000010010","000000000000000001","000000000000001101","000000000000000000","000000000000010110","000000000000000000","000000000000101000","000000000000000001","000000000000010110","000000000000001010","000000000000000000","000000000000000011","111111111111110011","000000000000010000","000000000000011010","000000000000000000","000000000000001000","111111111111111111","000000000000011100","000000000000000000","111111111111011101","000000000000011001","111111111111110100","000000000000000100","000000000000001011","000000000000001110","000000000000010010","000000000000011011","000000000000000110","000000000000010000","000000000000000000","111111111111111001","000000000000010011","111111111111111011","111111111111111000","000000000000001000","000000000000100100","000000000000010110","000000000000001101","000000000000001110","111111111111100001","111111111111011111","111111111111111100","111111111111111001","000000000000011000","000000000000001101","000000000000010011","000000000000111011","000000000000001100","000000000000000110","000000000000001000","000000000000000010","000000000000010001","000000000000001100","111111111111110110","000000000000100100","000000000000100010","111111111111101111","000000000000001001","000000000000000101","111111111111110101","111111111111111111","000000000000100001","000000000000010010","000000000000010010","000000000000000011","111111111111100100","000000000000010100","000000000000000100","000000000000000111","000000000000010111","000000000000010001","000000000000010011","000000000000000110","000000000000001100","000000000000000100","111111111111101001","111111111111111010","111111111111111010","000000000000001100","111111111111110001","111111111111100111","000000000000001110","000000000000000000","000000000000000111","000000000000000011","111111111111011011","000000000000010001","000000000000011011","000000000000000010","111111111111111010","000000000000011110","000000000000010100","111111111111110011","111111111111111010","111111111111110100","111111111111110000","000000000000010011","111111111111111111","111111111111100110","111111111111111001","111111111111111010","111111111111101000","000000000000000111","000000000000001011","000000000000001100","000000000000000101","111111111111100111","000000000000010111","111111111111101001","000000000000010010","111111111111111110","000000000000000111","000000000000011000","000000000000100100","111111111111110011","000000000000011001","111111111111001110","111111111111011100","000000000000011101","000000000000101011","000000000000001010"),
("000000000000010101","111111111111101011","000000000000000001","111111111111111101","111111111111100101","000000000000001110","000000000000000010","111111111111110000","111111111111101100","000000000000011000","000000000000000111","000000000000000001","000000000000110111","000000000000010000","000000000000000000","000000000000101011","111111111111101010","000000000000000000","111111111111101001","000000000000011101","111111111111111101","111111111111011010","111111111111110110","111111111111111100","111111111111111011","000000000000000101","111111111111001001","000000000000111000","111111111111100100","000000000000101000","000000000000011001","000000000000010000","000000000000100010","000000000000011011","000000000000000000","000000000000000011","000000000000000010","000000000000011001","111111111111110101","111111111111110010","000000000000000110","000000000000001000","000000000000010111","000000000000001000","000000000000010010","000000000000011010","000000000000000101","111111111111101010","000000000000000000","111111111111010010","111111111111101011","111111111111110000","000000000000000010","000000000000110000","000000000000010100","000000000000001011","000000000000010100","000000000000001010","000000000000001001","000000000000000111","000000000000001011","000000000000101010","000000000000001010","000000000000001101","000000000000100100","000000000000000111","111111111111111011","000000000000001110","000000000000010110","111111111111100101","000000000000000011","000000000000001010","111111111111101100","000000000000001001","000000000000010001","000000000000001000","000000000000010000","000000000000100100","000000000000000000","111111111111101101","000000000000010111","000000000000011101","111111111111101101","111111111111011100","000000000000001111","111111111111111100","111111111111111011","111111111111101101","111111111111111111","000000000000010011","000000000000010001","000000000000010000","111111111110111111","000000000000011100","000000000000000101","000000000000100101","111111111111101100","000000000000010011","000000000000100100","000000000000001110","111111111111111111","111111111111011111","000000000000001000","000000000000001010","111111111111100101","111111111111110111","000000000000010010","000000000000001110","111111111111100101","111111111111110010","111111111111111011","000000000000001100","000000000000001110","111111111111111111","111111111111110000","111111111111101010","000000000000011000","000000000000010011","000000000000001011","000000000000101100","000000000000101110","111111111111100101","000000000000010000","111111111111101111","111111111111011011","000000000000100010","000000000000100110","000000000000011111"),
("000000000000011110","111111111111111100","000000000000000000","000000000000001111","000000000000101000","111111111111110101","000000000000011110","111111111111111010","111111111111110001","111111111111100111","111111111111110001","000000000000000011","000000000000010100","000000000000001101","111111111111110101","111111111111111111","111111111111011110","000000000000011110","111111111111111111","111111111111101110","111111111111111100","111111111111010010","111111111111011011","000000000000010010","000000000000011100","000000000000001110","111111111111001010","000000000000101000","111111111111010001","000000000000001001","111111111111111100","000000000000011111","000000000000001000","000000000000100101","111111111111101111","111111111111101111","000000000000001011","111111111111111111","111111111111011010","111111111111101011","000000000000001101","000000000000001101","000000000000000001","000000000000011110","000000000000000100","000000000000010000","111111111111110011","111111111111110001","000000000000001010","000000000000000000","111111111111101111","111111111111111000","000000000000001001","000000000000010011","000000000000001001","111111111111110011","000000000000000011","000000000000001100","000000000000001111","000000000000000001","000000000000010100","000000000000011000","000000000000101010","000000000000010010","000000000000000001","000000000000011100","000000000000011000","111111111111110101","000000000000101011","111111111111100101","000000000000001010","000000000000001011","111111111111010001","000000000000101001","000000000000000100","111111111111110100","111111111111111001","000000000000100010","000000000000010000","111111111111101011","000000000000001111","000000000000011011","111111111111010111","111111111111101001","000000000000001101","000000000000001000","111111111111111100","000000000000000000","000000000000001011","000000000000001001","111111111111111011","000000000000000011","111111111110110011","000000000000100000","000000000000011101","000000000000100111","000000000000000000","000000000000011000","000000000000001110","000000000000010000","111111111111101110","000000000000001100","000000000000011110","111111111111110111","111111111111011010","000000000000000000","000000000000001000","000000000000101010","111111111111010101","111111111111100101","000000000000000000","111111111111111000","111111111111110001","111111111111110001","000000000000001101","000000000000011000","000000000000010100","000000000000000100","000000000000000111","000000000000001010","000000000000010000","111111111111011100","000000000000011010","111111111111100001","111111111111010100","000000000000101111","000000000000011110","000000000000011011"),
("000000000000011110","111111111111010100","000000000000010011","000000000000011110","000000000001011000","111111111111110000","000000000000011101","111111111111110010","111111111111111100","111111111111111001","111111111111110111","000000000000001101","111111111111110111","000000000000001010","111111111111111000","000000000000011011","111111111111110100","000000000000011101","000000000000000000","111111111111111100","000000000000001100","111111111111100010","111111111111110001","111111111111111101","000000000000001011","000000000000001100","111111111111011000","000000000000011100","111111111111100100","000000000000011001","000000000000001011","111111111111111101","000000000000011011","000000000000011001","111111111111100100","000000000000000010","000000000000000110","111111111111110111","111111111111101100","111111111111101110","000000000000010010","111111111111111111","111111111111111001","000000000000000000","000000000000001001","000000000000000000","111111111111011001","111111111111011000","111111111111101100","111111111111111100","111111111111111110","000000000000001000","000000000000011100","000000000000100011","000000000000010001","000000000000000011","000000000000001100","111111111111111011","000000000000010000","111111111111101011","000000000000011111","000000000000100001","000000000000001000","111111111111101111","000000000000011101","000000000000100001","000000000000010111","111111111111101001","000000000000001000","111111111111000111","111111111111111100","000000000000010011","111111111111101110","000000000000010110","111111111111110000","111111111111111110","000000000000010111","000000000000110001","000000000000000111","111111111111101010","111111111111101011","000000000000011000","111111111111011010","000000000000001000","111111111111110011","111111111111110000","111111111111111001","000000000000001001","111111111111100011","000000000000011001","111111111111001111","111111111111111110","111111111110110001","000000000000100111","000000000000010100","000000000000110000","111111111111111001","000000000000010011","111111111111110111","000000000000000000","111111111111101001","000000000000010010","000000000000110000","111111111111111010","111111111111110011","000000000000000101","000000000000011010","000000000000000100","111111111111111010","000000000000010011","000000000000000010","000000000000001110","111111111111101010","000000000000000011","111111111111110111","000000000000010110","111111111111111001","000000000000001000","000000000000001100","000000000000100111","000000000000111000","000000000000001000","000000000000000010","000000000000000000","111111111111101110","000000000000100101","000000000000100110","000000000000000100"),
("000000000000000111","111111111111111110","000000000000010111","000000000000001000","000000000001100010","111111111111100101","000000000000000101","111111111111100010","000000000000001011","111111111111110011","111111111111101011","111111111111111110","111111111111111101","000000000000011001","000000000000001100","000000000000011101","111111111111110101","000000000000010111","000000000000000100","111111111111111000","000000000000000010","111111111111110001","000000000000101001","000000000000010000","000000000000001010","000000000000000111","111111111111110001","000000000000010000","000000000000000110","000000000000010110","111111111111110010","000000000000000000","111111111111110100","000000000000000100","111111111111111000","111111111111101110","000000000000100001","000000000000001000","111111111111111011","111111111111111110","000000000000001110","000000000000010000","111111111111011011","000000000000001100","111111111111111010","000000000000001100","111111111111110010","111111111111011011","000000000000011110","000000000000011010","111111111111101010","111111111111110001","000000000000001011","111111111111101110","000000000000010101","000000000000001100","000000000000001000","000000000000010001","000000000000001110","000000000000001100","000000000000100101","000000000000011111","000000000000010100","111111111111110110","111111111111111110","000000000000011101","111111111111111110","111111111111110000","000000000000010110","111111111111011000","111111111111101100","000000000000010011","000000000000000001","000000000000011110","111111111111101101","111111111111111000","000000000000010001","000000000000010101","000000000000000111","111111111111101011","000000000000001110","111111111111111100","111111111111111100","000000000000100011","000000000000000010","000000000000010011","111111111111111011","111111111111111011","111111111111111100","111111111111110110","111111111111011011","000000000000011001","111111111110101011","000000000000010011","000000000000001011","000000000000100001","000000000000000011","111111111111110101","111111111111110111","111111111111011001","000000000000000110","111111111111110110","000000000000001111","000000000000001011","111111111111111101","111111111111111101","000000000000001110","000000000000000101","111111111111111110","111111111111111010","000000000000010011","000000000000001000","111111111111110100","000000000000000101","111111111111100100","000000000000111101","111111111111101001","000000000000001001","000000000000000010","000000000000011110","000000000000100110","000000000000001110","111111111111110001","111111111111111111","111111111111110110","111111111111111100","000000000000101011","000000000000010100"),
("000000000000001111","000000000000001001","000000000000001011","000000000000001101","000000000000101110","111111111111100010","000000000000000100","111111111111110011","111111111111111001","111111111111110001","111111111111111001","000000000000100001","000000000000000001","000000000000000000","111111111111110000","000000000000000000","000000000000000000","000000000000101000","000000000000011100","000000000000010101","000000000000001011","000000000000001110","000000000000011011","000000000000000000","000000000000010001","111111111111101001","111111111111110010","000000000000010110","000000000000011001","000000000000001111","111111111111111101","111111111111100000","000000000000001011","000000000000011111","000000000000000011","111111111111110100","000000000000000000","111111111111100101","000000000000000000","000000000000001101","000000000000011100","111111111111110101","111111111110110010","111111111111111010","111111111111110111","111111111111101010","111111111111100000","111111111111011100","000000000000010110","000000000000010010","000000000000000111","111111111111111010","000000000000101000","000000000000000010","111111111111111101","111111111111110110","000000000000011000","000000000000001101","000000000000010100","000000000000010000","000000000000010000","000000000000010011","000000000000001111","000000000000010111","111111111111111111","000000000000100010","000000000000011010","111111111111100110","111111111111111101","111111111111111001","111111111111110010","000000000000011000","000000000000010000","111111111111111110","111111111111111100","000000000000001101","111111111111110011","000000000000100010","000000000000000111","111111111111111111","111111111111110110","000000000000010001","111111111111101111","000000000000010111","000000000000010001","111111111111110101","000000000000001011","111111111111111010","111111111111110000","111111111111101000","111111111111011011","000000000000000100","111111111110100111","000000000000000000","000000000000011001","000000000000000001","111111111111010011","000000000000001000","111111111111100010","111111111111100100","111111111111110101","000000000000010010","000000000000101110","111111111111111100","111111111111111110","111111111111111111","111111111111111111","000000000000011001","000000000000000011","000000000000000000","000000000000100000","111111111111111100","111111111111110101","111111111111111101","111111111111110101","000000000000110100","000000000000000011","000000000000000001","111111111111101110","111111111111111001","000000000000110000","000000000000010100","111111111111111010","000000000000011110","111111111111110010","111111111111111100","000000000000110010","111111111111111000"),
("000000000000010011","111111111111111111","000000000000011100","000000000000100001","000000000000000000","000000000000000000","000000000000010000","000000000000000000","000000000000001001","111111111111110000","000000000000000001","000000000000100001","111111111111100101","000000000000011010","111111111111101000","000000000000010101","000000000000101010","000000000000001011","000000000000011001","111111111111111111","000000000000010100","000000000000001111","000000000000101110","000000000000000111","000000000000001011","111111111111101110","111111111111100100","111111111111110010","000000000000111010","000000000000010100","111111111111100111","111111111111100110","111111111111110100","000000000000011001","000000000000000000","000000000000000101","000000000000000100","111111111111101101","111111111111101111","000000000000000000","000000000000000010","111111111111101111","111111111110101010","111111111111110111","111111111111111010","111111111111111010","111111111111110110","111111111111111111","000000000000011011","000000000000011110","111111111111101101","000000000000000000","000000000000011110","111111111111100111","111111111111111101","000000000000011010","000000000000001000","000000000000100000","111111111111111111","000000000000000001","000000000000100100","000000000000001011","000000000000100100","000000000000001001","111111111111011111","000000000000001111","000000000000001001","111111111111110111","000000000000000110","000000000000010001","000000000000001011","000000000000100001","000000000000000000","111111111111000110","111111111111111100","111111111111111000","000000000000001111","000000000000000110","111111111111101111","111111111111111100","000000000000000011","000000000000001000","000000000000000000","000000000000110110","000000000000001011","111111111111110110","111111111111110110","000000000000000000","000000000000000000","111111111111100001","111111111111011010","000000000000001100","111111111110101001","111111111111110000","000000000000001110","111111111111111110","111111111111101000","111111111111101100","111111111111001101","000000000000100101","111111111111101100","111111111111111010","000000000000100101","000000000000000010","000000000000001101","111111111111111110","000000000000000011","000000000000000110","000000000000010111","111111111111111000","000000000000001011","111111111111111100","111111111111101000","000000000000001100","000000000000000100","000000000000110011","111111111111110101","111111111111111001","111111111111110101","111111111111110011","000000000001000001","111111111111111110","000000000000000100","000000000000001100","111111111111011101","111111111111111011","000000000000011000","000000000000001011"),
("000000000000011111","000000000000000000","000000000000001011","000000000000010001","000000000000001100","000000000000001000","000000000000000011","000000000000011000","111111111111101011","000000000000000010","111111111111111110","000000000000000111","000000000000000111","000000000000011101","000000000000001100","000000000000001010","000000000000011011","000000000000011100","000000000000011010","000000000000010011","111111111111111001","000000000000000100","000000000000111111","000000000000001000","000000000000000011","111111111111101110","111111111111111111","111111111111100100","000000000000010111","000000000000011100","111111111111111000","111111111111011110","111111111111110011","000000000000011000","000000000000001000","000000000000001101","000000000000100011","000000000000000010","111111111111110101","000000000000001011","000000000000010111","111111111111111011","111111111110111110","111111111111011111","111111111111110010","111111111111100111","111111111111111011","111111111111110101","000000000000001000","111111111111111111","111111111111111101","000000000000000001","111111111111111000","000000000000010010","000000000000001110","000000000000100100","000000000000010111","000000000000001110","111111111111111001","111111111111110110","000000000000000100","111111111111111101","000000000000000001","000000000000000101","111111111111011101","000000000000011001","000000000000001011","111111111111101101","111111111111111010","111111111111111101","000000000000001100","000000000000011000","000000000000000000","111111111110111111","111111111111110110","000000000000010000","000000000000001001","000000000000010011","000000000000001000","111111111111110100","000000000000000011","111111111111100110","000000000000000100","000000000000110001","111111111111110110","111111111111101110","000000000000011101","111111111111111100","111111111111110000","111111111111000111","111111111111111100","000000000000010101","111111111110100011","111111111111100011","111111111111101100","000000000000010101","111111111110111000","111111111111011101","111111111111100010","000000000000101110","111111111111011011","000000000000001111","000000000000001101","111111111111101010","000000000000001001","111111111111101010","000000000000000000","111111111111110110","000000000000010100","111111111111111011","000000000000000100","000000000000000110","000000000000000000","000000000000000110","000000000000010110","000000000000100111","111111111111111011","000000000000000101","000000000000001011","111111111111111010","000000000000101111","000000000000010001","111111111111111000","000000000000010100","111111111111101011","111111111111111100","000000000000100011","000000000000000010"),
("000000000000101111","111111111111101111","000000000000001010","000000000000010001","111111111111110100","000000000000000111","000000000000001111","000000000000101000","000000000000000001","111111111111100010","000000000000010101","000000000000001000","111111111111110111","000000000000000011","000000000000001011","000000000000000011","000000000000001111","000000000000010111","000000000000100111","000000000000001110","000000000000001101","000000000000001000","000000000000011010","000000000000001110","000000000000011010","111111111111111101","111111111111111100","111111111111111000","111111111111100011","000000000000010010","111111111111111000","111111111111011001","000000000000000111","000000000000010101","000000000000011101","111111111111110001","000000000000100000","000000000000000100","000000000000001100","000000000000000011","000000000000001010","000000000000000010","111111111111101100","000000000000000100","111111111111110100","111111111111010111","111111111111111000","111111111111100011","000000000000000111","111111111111101110","111111111111110101","111111111111110100","000000000000000100","111111111111111000","000000000000001000","000000000000010010","111111111111111011","111111111111110110","000000000000000000","111111111111111101","000000000000010010","000000000000000011","000000000000000000","000000000000010110","000000000000000101","000000000000011010","000000000000001000","111111111111100111","000000000000000000","000000000000000011","000000000000000000","000000000000011000","000000000000000100","111111111110111011","111111111111111111","111111111111110001","000000000000000011","000000000000010111","000000000000001010","111111111111111100","000000000000001110","111111111111110101","000000000000010001","000000000000011101","000000000000000110","000000000000000010","000000000000001010","000000000000001001","000000000000000000","111111111111000111","111111111111111101","000000000000001110","111111111110110000","000000000000000100","111111111111101001","111111111111111110","111111111111010110","111111111111110000","111111111111010101","000000000000010100","111111111111110110","000000000000100111","000000000000001100","111111111111100111","111111111111110110","000000000000000110","000000000000001100","111111111111111111","111111111111110100","000000000000011011","000000000000001110","000000000000000111","111111111111110001","111111111111100110","000000000000010000","000000000000010101","000000000000000100","000000000000000000","000000000000000111","111111111111101010","000000000000101000","000000000000001111","000000000000010111","000000000000000111","111111111111101000","111111111111100001","000000000000110110","000000000000001001"),
("000000000000111101","111111111111110001","111111111111111100","000000000000001101","111111111111111000","111111111111111101","111111111111111100","000000000000100101","111111111111111000","000000000000000000","000000000000010000","000000000000000010","000000000000001000","111111111111111111","111111111111101110","000000000000001011","000000000000001001","000000000000010001","000000000000100111","000000000000000100","000000000000010010","000000000000101001","000000000000010110","000000000000000111","000000000000010110","000000000000001000","000000000000000110","111111111111010110","111111111110111110","000000000000100101","111111111111111111","111111111111100111","111111111111110111","000000000000011100","000000000000001011","111111111111100100","000000000000001001","111111111111110011","000000000000001101","111111111111110111","111111111111111110","111111111111111101","111111111111011100","111111111111111000","111111111111111011","111111111111111110","111111111111110001","111111111111101101","000000000000000100","111111111111101000","000000000000001101","000000000000011111","111111111111110111","111111111111010100","000000000000000111","000000000000100001","000000000000000000","000000000000000000","000000000000001110","111111111111101100","000000000000001111","000000000000100000","111111111111101101","000000000000010011","111111111111010111","111111111111111111","000000000000000111","000000000000000001","111111111111101010","111111111111111101","111111111111101000","000000000000010001","000000000000010101","111111111111001001","111111111111110000","111111111111110101","000000000000100010","000000000000001100","111111111111111110","000000000000010100","000000000000000111","111111111111111000","000000000000001001","000000000000000011","000000000000000101","111111111111110000","000000000000010110","111111111111110001","111111111111111110","111111111111010110","111111111111110001","000000000000000001","111111111111000010","111111111111110101","111111111111101100","111111111111110101","111111111111010110","111111111111101000","111111111111110000","000000000000101001","000000000000000100","000000000000100000","000000000000010001","000000000000010000","000000000000000100","000000000000010100","000000000000000111","111111111111111010","111111111111110110","000000000000011000","111111111111110010","111111111111110001","000000000000001101","000000000000000000","000000000000100100","000000000000000001","111111111111111000","111111111111101101","000000000000000010","111111111111111101","000000000000100000","000000000000001101","111111111111110101","000000000000001110","111111111111110001","111111111111101101","000000000000100011","111111111111111100"),
("000000000000101001","111111111111110011","000000000000000000","000000000000000011","111111111111110000","000000000000000100","111111111111110001","000000000000100100","111111111111101100","111111111111110111","000000000000001111","000000000000000011","111111111111110101","111111111111111100","111111111111100110","000000000000010100","000000000000000000","000000000000001110","000000000000001110","000000000000000000","111111111111110110","000000000000101110","000000000000001010","000000000000010100","000000000000011001","111111111111100010","000000000000011011","111111111111001101","111111111111001101","111111111111111110","111111111111100111","111111111111101000","111111111111111000","111111111111111010","000000000000000011","111111111111111001","000000000000000001","000000000000001101","000000000000101100","000000000000000111","111111111111110011","111111111111111010","111111111111101101","111111111111010101","000000000000010100","111111111111011110","111111111111111101","111111111111101110","000000000000010101","000000000000000011","111111111111111001","000000000000010110","000000000000000101","111111111111010011","111111111111101100","111111111111111111","000000000000010010","000000000000000011","000000000000000010","111111111111111001","000000000000100000","111111111111110111","111111111110111011","000000000000011010","111111111111010100","000000000000001100","000000000000101110","111111111111111101","111111111111011011","111111111111110011","111111111111111110","000000000000010010","000000000000011100","111111111111000101","111111111111001011","111111111111100100","111111111111110110","111111111111110011","111111111111101010","000000000000001111","000000000000101101","111111111111110011","111111111111111010","000000000000011010","000000000000010101","111111111111100001","111111111111100100","000000000000001101","000000000000001101","111111111111100001","000000000000001111","000000000000011001","111111111111011001","111111111111101000","000000000000000000","111111111111100010","111111111111110010","111111111111000011","111111111111101111","000000000000011011","111111111111111101","000000000000000111","000000000000001100","000000000000010100","000000000000000001","000000000000011110","000000000000001000","111111111111100111","000000000000001000","000000000000001101","000000000000011101","000000000000000001","000000000000000110","000000000000000010","000000000000100110","111111111111110100","111111111111111000","111111111111011101","000000000000010011","111111111111101110","000000000000101100","111111111111110110","111111111111100010","111111111111111100","111111111111011110","111111111111010100","000000000000100010","111111111111110110"),
("000000000000010111","000000000000101101","000000000000010110","111111111111010001","111111111111011100","111111111111101100","111111111111111101","111111111111111001","111111111111010111","000000000000000100","111111111111110010","000000000000001011","111111111111001100","111111111111101011","111111111111101100","111111111111011010","000000000000000100","111111111111101001","000000000000010000","111111111111100011","111111111111011100","111111111111111001","111111111111101011","000000000000001011","000000000000010101","111111111111101111","000000000000000000","111111111111000101","111111111111101000","000000000000010000","000000000000000101","111111111111011001","000000000000010010","000000000000000010","000000000000000010","111111111111111000","000000000000010000","000000000000000011","000000000000100000","000000000000000000","000000000000011010","111111111111111100","111111111111001100","111111111111000011","000000000000011110","111111111111111001","111111111111110011","111111111111111101","000000000000011001","000000000000000001","000000000000001000","000000000000100100","111111111111110000","111111111111100110","111111111111110101","000000000000000010","000000000000011010","000000000000000010","000000000000000001","111111111111110010","000000000000010011","111111111111111011","111111111110111011","111111111111110100","111111111111100110","000000000000010001","000000000000000000","111111111111111111","111111111111110111","000000000000000101","111111111111101101","111111111111100101","000000000000001001","111111111111101110","111111111111100011","000000000000000111","000000000000001011","111111111111101000","000000000000001110","111111111111111101","000000000000010010","000000000000000101","000000000000001111","111111111111100101","111111111111100000","111111111111101110","111111111111110111","000000000000001000","000000000000010010","111111111111011010","000000000000010100","111111111111111011","111111111111011010","111111111111110001","111111111111111100","111111111111100110","111111111111011011","111111111111011010","111111111111110111","000000000000101001","000000000000011100","000000000000010010","111111111111101011","000000000000000011","111111111111111011","000000000000010000","000000000000000000","111111111111110101","111111111111111000","111111111111101110","111111111111111100","111111111111110100","000000000000011100","000000000000000011","000000000000000111","000000000000000100","000000000000011001","111111111111110100","111111111111111010","111111111111100001","000000000000000110","000000000000001010","111111111111011111","111111111111110011","111111111111111110","111111111111011111","111111111111111110","111111111111101011"),
("000000000000110011","000000000000001011","000000000000010101","111111111111110101","000000000000011100","000000000000001010","000000000000010011","111111111111010110","111111111111011011","111111111111101001","111111111111000111","000000000000011100","111111111111100011","111111111111100000","111111111111100110","111111111111100101","111111111111000100","111111111111111011","111111111111110010","111111111111011101","111111111111011111","000000000000011011","111111111111001111","111111111111110000","000000000000010110","000000000000000010","000000000000001010","111111111111100110","111111111111110010","000000000000001101","000000000000101000","111111111111011100","000000000000100010","000000000000000000","000000000000100001","000000000000000100","000000000000001100","000000000000011110","000000000000011010","000000000000001100","000000000000100010","000000000000001111","111111111111110001","111111111111110101","000000000000101111","111111111111100100","111111111111111010","000000000000010000","000000000000010101","000000000000010010","111111111111100000","000000000000011000","111111111111100000","000000000000001000","000000000000001011","000000000000000000","000000000000100010","111111111111011001","111111111111111011","000000000000010001","111111111111111100","111111111111001101","111111111111010001","000000000000000001","000000000000001010","000000000000010010","111111111111110111","111111111111110101","111111111111100111","000000000000000011","000000000000000001","111111111111111001","111111111111110110","111111111111110011","111111111111101111","000000000000000111","000000000000100000","111111111111010111","111111111111111101","000000000000001101","000000000000011101","000000000000100101","111111111111111111","111111111111100001","111111111111110001","111111111111110100","000000000000101111","111111111111111000","111111111111100111","111111111111100010","000000000000011011","111111111111101010","111111111111111011","111111111111110000","111111111111101111","111111111111100111","000000000000000000","000000000000100111","000000000000000001","000000000000001011","000000000000101100","000000000000000010","111111111111101001","000000000000001100","111111111111111111","000000000000000110","111111111111101101","111111111111011001","000000000000001010","111111111111111111","111111111111110000","000000000000000110","000000000000011011","111111111111111100","000000000000011001","111111111111100111","000000000000010001","000000000000101010","000000000000000011","000000000000011110","000000000000001101","000000000000101000","000000000000000011","111111111110111110","111111111111110010","111111111111100101","000000000000001110","111111111111110110"),
("000000000000011000","000000000000000110","000000000000101110","111111111111111011","000000000000010110","000000000000001100","111111111111101000","111111111111101101","000000000000001111","111111111111110111","111111111111011001","111111111111111101","111111111111111001","111111111111110111","000000000000000000","000000000000000000","111111111111100100","000000000000001001","000000000000010011","111111111111101110","111111111111111000","111111111111100110","111111111111001010","111111111111011111","111111111111111100","000000000000001000","000000000000001111","111111111111110010","111111111111111110","000000000000011100","000000000000010110","111111111111110110","111111111111110001","111111111111111111","000000000000010010","000000000000001101","000000000000001001","000000000000100111","000000000000010011","000000000000000101","000000000000100001","000000000000010110","000000000000001111","000000000000000000","000000000001000100","000000000000000110","000000000000010001","111111111111110000","000000000000011011","111111111111110100","111111111111100011","000000000000001000","111111111111100111","000000000000011001","111111111111111011","000000000000001100","000000000000000110","111111111111011101","111111111111101111","111111111111101101","111111111111110000","111111111111100010","111111111111100010","000000000000000100","111111111111101000","000000000000000010","111111111111111011","111111111111110011","111111111111111010","000000000000101110","111111111111101001","111111111111111101","111111111111111001","111111111111110000","111111111111111110","111111111111110111","000000000000010110","000000000000000000","111111111111110011","111111111111101111","000000000000100111","000000000000011001","000000000000010110","000000000000010010","111111111111110010","000000000000000010","000000000000100110","000000000000110001","111111111111111111","111111111111100110","000000000000100110","111111111111100110","111111111111111101","111111111111011011","111111111111101111","000000000000001101","000000000000000010","111111111111100110","000000000000000000","000000000000010110","000000000000011110","000000000000100001","111111111111011000","111111111111101101","111111111111111111","111111111111111000","111111111111101100","111111111111111010","000000000000001000","111111111111101100","111111111111100110","000000000000000001","000000000000011110","111111111111111001","000000000000010110","111111111111100111","111111111111111101","000000000000011001","000000000000001010","000000000000110001","000000000000001110","000000000000100101","000000000000000000","111111111111011001","111111111111110111","111111111111111110","111111111111111011","000000000000001000"),
("000000000000110010","000000000000001001","000000000000000101","111111111111110110","000000000000100101","000000000000011100","000000000000010101","000000000000000001","111111111111111011","111111111111101001","111111111111111110","000000000000101000","000000000000011100","111111111111100001","111111111111110011","000000000000010111","000000000000001011","111111111111111010","111111111111101101","000000000000000000","111111111111110100","000000000000000110","111111111111100011","111111111111111110","111111111111101111","000000000000001001","000000000000000011","111111111111110110","000000000000000011","000000000000000001","111111111111110111","000000000000001011","111111111111101001","111111111111111010","000000000000011001","111111111111111010","111111111111101101","111111111111110111","111111111111110010","111111111111101101","000000000000011011","000000000000010100","000000000000010111","000000000000010001","000000000000001011","111111111111100101","000000000000011111","000000000000000011","000000000000011000","000000000000011011","111111111111110111","111111111111101010","111111111111101101","000000000000011011","111111111111101100","111111111111011101","000000000000011011","111111111111100100","000000000000000000","000000000000001001","000000000000001000","111111111111111101","111111111111111101","111111111111110010","111111111111101000","111111111111110010","111111111111101000","000000000000011000","111111111111110101","000000000000011001","000000000000010011","111111111111101100","000000000000000000","111111111111111001","111111111111110010","000000000000010011","111111111111110110","111111111111101010","111111111111111011","111111111111110111","111111111111111111","111111111111111100","000000000000010110","000000000000001110","000000000000001001","111111111111000011","000000000000011000","111111111111111001","000000000000001001","111111111111100101","111111111111111101","000000000000001101","000000000000011101","111111111111000111","000000000000010010","000000000000010101","111111111111100111","000000000000000000","000000000000001100","000000000000100010","000000000000011111","000000000000000010","000000000000001100","000000000000000000","000000000000000000","000000000000000111","000000000000000010","111111111111111001","111111111111100000","111111111111111000","000000000000001001","000000000000000010","000000000000100101","111111111111110001","111111111111110011","000000000000001000","000000000000100001","000000000000101111","000000000000000001","000000000000011000","111111111111110100","111111111111100110","000000000000000001","111111111111101001","111111111111111000","111111111111111010","000000000000011111","000000000000001110"),
("111111111111101001","111111111111110101","111111111111100010","000000000000000001","000000000000011101","111111111111100010","000000000000100000","000000000000000010","111111111111101101","000000000000011100","000000000000100011","000000000000001111","111111111111010001","111111111111100010","111111111111100010","111111111111111010","000000000000010100","000000000000101001","111111111111100001","000000000000011100","111111111111100110","000000000000010010","000000000000001011","000000000000010011","000000000000101011","111111111111010111","000000000000001101","111111111111110101","111111111111110000","000000000000010000","111111111111010111","111111111111111111","000000000000001110","000000000000010010","000000000000000110","000000000000001001","111111111111111000","111111111111011000","111111111111101111","111111111111011100","000000000000000101","111111111111111001","111111111111111010","000000000000011001","111111111111111110","111111111111010110","111111111111110011","111111111111111101","111111111111111111","111111111111111100","000000000000100101","000000000000100000","000000000000011110","000000000000000111","111111111111011100","111111111111101010","111111111111110000","000000000000001111","000000000000001001","000000000000001110","000000000000000101","111111111111101111","000000000000100111","000000000000011111","000000000000001101","000000000000101110","000000000000101000","111111111111111110","111111111111110101","000000000000110010","111111111111101011","111111111111101110","000000000000000100","000000000000001000","111111111111110110","000000000000001111","111111111111010101","000000000000001001","111111111111101010","000000000000011011","000000000000011011","111111111111101101","000000000000000001","111111111111101001","000000000000001110","000000000000101000","111111111111111000","000000000000000100","111111111111110000","000000000000000011","111111111111110111","111111111111101110","000000000000010110","000000000000100111","111111111111110110","111111111111110100","000000000000010011","111111111111011011","000000000000001010","111111111111100111","000000000000010100","000000000000010001","000000000000011101","111111111111111101","000000000000001110","000000000000011110","111111111111110011","111111111111010100","000000000000000011","000000000000001101","111111111111101000","111111111111110101","000000000000101010","111111111111101100","111111111111100011","000000000000001000","000000000000000000","111111111111110010","000000000000001000","111111111111110110","000000000000001111","000000000000001010","111111111111111010","111111111111011010","000000000000011010","111111111111111100","000000000000010010","111111111111011111"),
("111111111111111000","111111111111111001","000000000000010101","000000000000001100","111111111111100111","111111111111111111","000000000000001001","111111111111010101","000000000000100011","000000000000001111","000000000000011101","111111111111101101","000000000000001110","111111111111111110","111111111111111101","000000000000011110","000000000000010110","000000000000001001","000000000000001111","000000000000000010","000000000000011110","000000000000000100","111111111111110010","111111111111001110","000000000000000000","111111111111100111","111111111111101100","000000000000000011","000000000000001111","000000000000000110","111111111111111010","111111111111111011","000000000000001110","111111111111111000","000000000000100000","111111111111001111","000000000000010110","000000000000011010","111111111111111001","111111111111111111","000000000000010000","000000000000011011","000000000000011111","111111111111101010","111111111111110111","000000000000011001","000000000000100011","000000000000001000","000000000000000001","111111111111111100","000000000000011010","111111111111111101","000000000000011101","111111111111111001","000000000000011100","000000000000010001","111111111111110001","000000000000011111","111111111111111101","000000000000001101","000000000000001000","000000000000000010","000000000000010100","111111111111011001","111111111111011000","000000000000001110","111111111111100111","111111111111100111","111111111111110000","000000000000100001","111111111111110110","000000000000010110","000000000000000100","000000000000010001","111111111111101011","111111111111111110","111111111111111100","111111111111110001","000000000000001010","000000000000000100","111111111111100010","111111111111111010","000000000000000000","000000000000001011","000000000000000100","000000000000011011","000000000000010001","111111111111111110","111111111111101001","000000000000011100","111111111111110111","000000000000000101","000000000000110101","000000000000001101","111111111111111110","000000000000001011","000000000000010010","000000000000000111","111111111111110011","000000000000000101","111111111111101100","000000000000001000","111111111111110101","111111111111111000","000000000000000101","111111111111101010","111111111111110000","000000000000010110","111111111111101100","000000000000010111","000000000000000100","000000000000000111","111111111111101101","000000000000000111","000000000000111011","000000000000001110","000000000000000000","000000000000010111","111111111111100111","000000000000010001","000000000000000111","111111111111111001","000000000000010110","000000000000110110","000000000000001011","111111111111011110","000000000000011001","111111111111010110"),
("111111111111111110","000000000000000001","000000000000011100","111111111111011010","000000000000010000","111111111111111011","111111111111111010","111111111111101011","111111111111110111","111111111111110000","111111111111101001","111111111111111100","000000000000000101","111111111111111101","000000000000100110","000000000000001100","000000000000011110","000000000000010010","000000000000001000","000000000000101001","111111111111101100","000000000000100011","000000000000010101","111111111111110011","000000000000001100","111111111111100100","000000000000010110","111111111111100110","000000000000010000","111111111111111010","111111111111111011","111111111111010100","111111111111011000","111111111111010111","111111111111110101","111111111111101110","000000000000011100","111111111111101010","111111111111111011","000000000000000101","111111111111100101","000000000000000000","000000000000000011","111111111111011111","000000000000010011","000000000000000000","000000000000000100","111111111111111010","000000000000101100","111111111111110001","111111111111101101","000000000000010001","111111111111110111","111111111111011001","000000000000000111","000000000000011101","111111111111111110","000000000000000000","000000000000011110","000000000000001010","111111111111101010","000000000000001001","000000000000000000","000000000000010100","111111111111010000","000000000000011101","000000000000001000","000000000000000000","000000000000100000","000000000000100011","111111111111011000","111111111111111101","111111111111011011","111111111111110011","111111111111100010","111111111111110011","000000000000000000","000000000000001000","000000000000011001","000000000000011101","111111111111110111","111111111111101001","000000000000010111","000000000000001111","111111111111011101","000000000000110110","000000000000000010","000000000000010110","000000000000001110","000000000000001111","111111111111101000","111111111111111110","111111111111110000","000000000000010001","000000000000001101","000000000000000000","000000000000010101","000000000000000000","111111111111100111","000000000000000100","000000000000000110","000000000000000001","111111111111101101","111111111111101000","000000000000100001","111111111111101001","000000000000001000","111111111111111100","111111111111111111","000000000000101111","000000000000010000","111111111111110111","111111111111101110","000000000000011100","000000000000011000","111111111111110001","000000000000001100","111111111111111110","000000000000001000","111111111111111011","000000000000010110","000000000000000110","111111111111111000","000000000000001101","000000000000011111","111111111111101110","000000000000011011","000000000000000011"),
("111111111111110111","111111111111011011","000000000000010010","111111111111100100","000000000000011101","111111111111101000","111111111111111010","000000000000000000","000000000000100110","000000000000011011","111111111111110011","111111111111100111","111111111111111001","000000000000001111","000000000000011011","000000000000001001","000000000000100111","000000000000010111","000000000000011100","000000000000101011","000000000000010100","000000000000010110","000000000000100111","000000000000011000","111111111111100110","111111111111111010","000000000000100001","111111111111110010","000000000000100101","111111111111101011","111111111111011010","111111111111111101","111111111111110101","111111111111100001","000000000000000001","000000000000000100","111111111111101000","000000000000000100","111111111111110001","000000000000011000","111111111111101010","111111111111111011","000000000000011001","000000000000000100","000000000000001000","000000000000010100","000000000000001010","111111111111010110","000000000000100110","111111111111111000","000000000000110100","000000000000000000","111111111111111101","111111111111110011","000000000000010111","000000000000000010","111111111111011000","000000000000001010","000000000000010000","000000000000001111","000000000000000100","111111111111111111","000000000000000010","000000000000000010","111111111111111101","000000000000000000","000000000000001001","000000000000000101","000000000000001011","111111111111110000","000000000000001011","000000000000011110","000000000000000000","000000000000010101","111111111111100110","111111111111101011","111111111111101100","111111111111100110","000000000000010100","000000000000011100","111111111111100011","111111111111011000","000000000000001110","000000000000100111","111111111111110111","111111111111111111","000000000000011010","111111111111111101","111111111111101110","111111111111111111","111111111111101010","111111111111101011","111111111111110111","000000000000010011","111111111111111001","111111111111110000","000000000000000101","111111111111111000","000000000000001111","000000000000000000","111111111111101110","111111111111110011","000000000000000001","000000000000010100","000000000000010010","000000000000001000","000000000000011000","000000000000001111","000000000000010000","000000000000000010","111111111111111011","111111111111110010","000000000000000011","000000000000101001","000000000000100110","000000000000001000","000000000000001000","000000000000001000","111111111111110001","000000000000010010","111111111111111110","111111111111110100","111111111111101100","000000000000001110","111111111111110110","111111111111011100","000000000000000101","000000000000001111"),
("111111111111011011","000000000000001011","000000000000001001","000000000000001101","000000000000101010","111111111111101100","111111111111111010","000000000000000101","000000000000110011","000000000000011100","000000000000010011","111111111111101001","000000000000100010","000000000000000111","000000000000100011","111111111111111001","000000000000100111","111111111111110000","000000000000001101","000000000000101100","000000000000000101","000000000000100001","000000000000001011","111111111111100110","111111111111101100","000000000000011100","000000000000001101","111111111111111111","000000000000010110","111111111111101111","111111111111100000","000000000000010000","111111111111101110","111111111111010001","111111111111101011","000000000000100011","111111111111111111","000000000000011001","111111111111110000","111111111111111111","111111111111010001","111111111111101000","000000000000011001","111111111111111011","111111111111110110","000000000000011111","000000000000101011","111111111110101010","000000000000010100","111111111111110110","000000000000011010","111111111111111111","111111111111110010","111111111111010110","000000000000000000","000000000000100100","111111111111001110","111111111111110101","000000000000000111","000000000000000001","111111111111101011","111111111111110011","000000000000000000","000000000000000110","000000000000001001","111111111111100111","111111111111111111","111111111111110110","000000000000010000","111111111111111100","000000000000001111","000000000000010000","000000000000001101","000000000000100000","000000000000000110","000000000000011010","111111111111111100","000000000000001110","000000000000100010","000000000000010010","111111111111110000","000000000000000000","000000000000001001","111111111111110111","000000000000000011","000000000000010000","000000000000000110","000000000000000001","111111111111110110","000000000000001111","111111111111111000","111111111111011110","000000000000001101","111111111111111101","111111111111111000","111111111111011100","000000000000001000","000000000000011100","000000000000001001","111111111111011011","111111111111110100","111111111111100111","000000000000001000","000000000000001101","000000000000010110","000000000000011000","111111111111111001","000000000000001101","111111111111111011","111111111111110111","111111111111110101","000000000000000011","000000000000011100","000000000000001110","000000000000010101","111111111111111110","000000000000000101","111111111111110110","111111111111101100","000000000000000110","000000000000000000","111111111111101001","111111111111111110","000000000000100110","000000000000000000","111111111110111000","111111111111111101","111111111111101001"),
("111111111111010000","111111111111111001","000000000000000110","111111111111111010","000000000000100011","111111111111111101","111111111111101100","000000000000100101","000000000000011011","111111111111110001","111111111111110010","000000000000011100","000000000000001000","111111111111111100","000000000000100010","111111111111111100","000000000000011111","000000000000010110","000000000000100000","000000000000000000","000000000000000011","000000000000001110","111111111111111111","111111111111111110","000000000000000100","111111111111110010","000000000000010111","111111111111101101","000000000000001100","111111111111011111","111111111111101000","111111111111101101","000000000000001110","111111111111010100","000000000000000010","000000000000011010","000000000000000111","000000000000001011","111111111111100111","000000000000011100","111111111111110111","111111111111000110","000000000000100010","000000000000000100","000000000000010011","000000000000010010","000000000000000010","111111111111100111","000000000000011000","000000000000001000","000000000000011101","111111111111110101","111111111111111011","111111111111111011","111111111111110110","000000000000100011","111111111111100010","000000000000000001","000000000000001001","000000000000010000","111111111111101001","111111111111011100","111111111111111000","111111111111111011","111111111111010000","111111111111110000","111111111111011101","111111111111011010","000000000000011100","000000000000001010","111111111111110011","000000000000000111","000000000000001001","111111111111111000","000000000000010000","000000000000011101","000000000000010011","111111111111101010","111111111111111100","000000000000000011","111111111111101011","111111111111101110","111111111111111010","111111111111100100","111111111111110101","000000000000100100","000000000000011100","000000000000000111","111111111111110000","111111111111110111","111111111111100110","111111111111011110","000000000000010010","111111111111110000","000000000000000110","111111111111110001","111111111111111011","000000000000000101","111111111111100100","111111111111101111","111111111111011101","111111111111110100","111111111111110010","000000000000000010","000000000000010011","000000000000000111","000000000000001110","000000000000000001","000000000000000110","000000000000001100","000000000000010110","000000000000000101","000000000000001010","000000000000000001","000000000000011111","111111111111110011","111111111111101001","000000000000010011","111111111111101010","000000000000000001","111111111111110001","111111111111101111","111111111111100000","000000000000000101","000000000000010000","111111111111100001","000000000000011001","111111111111110100"),
("111111111111100011","111111111111111010","000000000000000110","111111111111110010","000000000000011000","111111111111101011","000000000000001000","000000000000010010","000000000000010011","000000000000000000","111111111111101010","000000000000001000","111111111111111111","000000000000000000","000000000000011111","111111111111110101","000000000000000110","111111111111111111","000000000000011101","000000000000000011","000000000000001111","000000000000100011","000000000000001000","111111111111111101","111111111111100101","111111111111110100","000000000000000011","111111111111110001","000000000000100000","111111111111110010","111111111111100101","111111111111101010","000000000000000010","111111111111100000","000000000000001111","111111111111111110","000000000000000011","000000000000000001","111111111111100101","111111111111111010","000000000000001100","111111111111010010","000000000000011011","111111111111111010","000000000000010000","111111111111110010","111111111111110011","111111111111111001","000000000000000111","111111111111111111","000000000000001111","111111111111110101","111111111111110010","000000000000001111","000000000000000001","000000000000001011","111111111111100110","111111111111111011","000000000000010100","000000000000000000","111111111111110010","111111111111100011","000000000000001110","111111111111101101","111111111110110010","000000000000011101","111111111111111000","111111111111110101","111111111111111001","000000000000001001","000000000000000100","111111111111101001","000000000000000101","000000000000010100","000000000000000000","111111111111111100","000000000000010101","111111111111110101","000000000000100010","000000000000001001","000000000000001011","111111111111101110","111111111111101100","111111111111000010","111111111111110010","000000000000010010","000000000000001011","000000000000000000","111111111111101000","111111111111111110","111111111111101110","111111111111111110","000000000000001001","111111111111100000","000000000000001110","111111111111011001","111111111111110101","000000000000001111","111111111111011111","000000000000000110","111111111111101010","000000000000010100","111111111111110010","111111111111111010","111111111111111100","111111111111110110","000000000000001111","000000000000000111","000000000000001011","000000000000001101","000000000000010100","111111111111111100","111111111111111100","111111111111111110","000000000000101110","111111111111011100","000000000000000001","000000000000000000","111111111111110001","111111111111101111","111111111111111011","111111111111101100","111111111111101100","000000000000011111","111111111111111110","111111111111110110","111111111111111111","000000000000001100"),
("111111111110111111","000000000000010010","111111111111111010","111111111111101101","000000000000101011","111111111111001110","111111111111111111","111111111111111000","000000000000000001","111111111111110010","000000000000000111","000000000000001100","000000000000001001","000000000000001100","000000000000000010","111111111111110010","111111111111101100","000000000000000001","000000000000100101","111111111111111100","000000000000001000","000000000000000010","000000000000001111","111111111111110001","111111111111101111","000000000000000110","000000000000000001","111111111111110001","000000000000010010","111111111111010011","111111111111100110","111111111111110110","111111111111111101","111111111111111000","000000000000100100","000000000000001100","111111111111111100","000000000000001010","111111111111110000","000000000000000111","111111111111111000","111111111111111000","111111111111111001","111111111111111101","000000000000000000","000000000000000010","111111111111111101","000000000000010001","000000000000010111","000000000000011100","000000000000010011","111111111111100000","111111111111110110","000000000000001000","000000000000001011","000000000000000000","111111111111111001","111111111111111110","000000000000000000","111111111111101101","111111111111111101","111111111111101010","111111111111101100","111111111111111110","111111111110110011","111111111111111100","111111111111100110","111111111111100000","000000000000001010","000000000000010001","000000000000001001","000000000000001100","111111111111111011","000000000000000011","111111111111111000","000000000000000000","111111111111101110","111111111111111001","000000000000001100","000000000000001000","111111111111110110","000000000000000000","111111111111100101","000000000000001000","000000000000001011","111111111111101010","000000000000010011","000000000000000000","111111111111111000","111111111111101100","111111111111111000","111111111111110010","000000000000001001","000000000000000010","000000000000000111","111111111111001010","111111111111110101","000000000000001100","111111111111110001","000000000000001111","111111111111100110","000000000000010011","111111111111100001","111111111111111101","111111111111110011","000000000000010011","000000000000000001","000000000000011101","111111111111110111","111111111111111001","000000000000001010","000000000000000110","111111111111111111","000000000000011100","000000000000110010","111111111111110100","111111111111110000","000000000000010110","111111111111110011","000000000000001011","000000000000011010","111111111111101101","000000000000001011","000000000000100111","000000000000000000","111111111111110101","000000000000010000","000000000000001101"),
("111111111111000010","000000000000010111","000000000000000000","111111111111110111","000000000000011001","111111111111101000","111111111111111000","111111111111111101","000000000000001111","000000000000000000","000000000000001101","000000000000011000","000000000000100000","111111111111111010","000000000000010100","000000000000001001","111111111111011100","000000000000010101","000000000000000010","000000000000010000","000000000000000100","111111111111111010","000000000000010001","111111111111100001","000000000000001100","111111111111111110","111111111111110100","000000000000011111","111111111111111110","111111111111010010","000000000000000100","000000000000001101","000000000000010110","111111111111110010","111111111111111101","000000000000010101","000000000000001001","111111111111101111","000000000000010100","000000000000001011","000000000000010111","111111111111110101","000000000000010001","111111111111110101","000000000000000111","000000000000000000","111111111111111010","000000000000001011","000000000000010110","000000000000010001","111111111111110110","111111111111100100","111111111111111001","000000000000010111","000000000000001110","000000000000011010","111111111111110110","000000000000001100","000000000000010110","111111111111101101","111111111111101010","111111111111111011","000000000000000101","000000000000000000","111111111111100100","000000000000100101","111111111111011011","111111111111111110","000000000000011001","000000000000010000","000000000000001100","111111111111110110","111111111111001011","111111111111110011","111111111111110011","000000000000010001","111111111111111111","000000000000010000","000000000000000110","000000000000000101","111111111111110001","111111111111110100","111111111111010011","111111111111111001","111111111111101101","000000000000000011","000000000000010011","111111111111110011","000000000000010001","111111111111111010","111111111111110111","111111111111110111","000000000000010110","111111111111111100","000000000000011000","000000000000000000","000000000000001111","000000000000010111","111111111111011000","111111111111110010","111111111111110101","000000000000010101","111111111111111011","111111111111101111","111111111111011010","000000000000001101","000000000000001011","000000000000011000","000000000000011001","000000000000000111","000000000000011101","000000000000001000","000000000000000000","000000000000001110","000000000000000000","111111111111010111","111111111111110111","111111111111110111","111111111111110101","000000000000010001","000000000000010001","111111111111110000","000000000000001011","000000000000011010","111111111111111001","000000000000100111","000000000000010111","111111111111111010"),
("111111111111001001","000000000000100011","000000000000010000","111111111111111010","000000000000101101","111111111111110111","111111111111111100","111111111111111110","000000000000001000","000000000000001010","111111111111101010","000000000000010100","000000000000000101","000000000000010010","000000000000011011","000000000000000100","111111111111111011","000000000000100011","000000000000000000","000000000000011001","111111111111110101","000000000000010010","000000000000001010","111111111111010100","000000000000010110","111111111111100010","000000000000001100","000000000000001000","111111111111110101","111111111111011010","000000000000001001","000000000000000001","000000000000010011","000000000000000100","000000000000010000","111111111111111111","000000000000000000","111111111111101001","000000000000010011","000000000000000000","000000000000000100","000000000000000000","000000000000011000","000000000000001011","111111111111101001","111111111111010101","000000000000000000","000000000000010100","000000000000000010","000000000000010011","000000000000000000","000000000000000010","000000000000011001","000000000000001001","000000000000010011","111111111111111001","111111111111111001","000000000000010000","000000000000001111","000000000000001000","111111111111100001","111111111111110000","111111111111111101","111111111111111110","111111111111110011","000000000000010011","111111111111011111","111111111111111011","000000000001000001","000000000000000000","000000000000000110","000000000000010000","111111111111000111","111111111111111101","111111111111110111","000000000000010100","000000000000000000","111111111111110010","111111111111111111","000000000000000010","000000000000000010","000000000000000100","000000000000000010","000000000000101101","111111111111110001","000000000000001000","111111111111110100","111111111111101000","000000000000010000","111111111111101110","000000000000001110","111111111111110011","000000000000000101","111111111111111110","000000000000000100","111111111111011101","111111111111011111","000000000000000111","111111111111001101","111111111111101101","111111111111110001","000000000000011101","111111111111110100","000000000000000101","111111111111110000","111111111111111111","000000000000011100","000000000000010010","000000000000010011","000000000000001101","000000000000010000","111111111111111001","111111111111110001","000000000000001001","000000000000011011","111111111111100100","111111111111111011","111111111111110010","111111111111111110","000000000000011110","000000000000011101","111111111111110101","000000000000000000","000000000000001010","111111111111110001","000000000000011111","000000000000011010","000000000000010001"),
("111111111111101011","000000000000010000","000000000000001100","000000000000000111","111111111111101010","000000000000000010","000000000000011011","000000000000000001","111111111111110101","000000000000001000","000000000000000001","000000000000001111","000000000000111111","111111111111101110","000000000000001110","000000000000101111","111111111111111010","000000000000010110","000000000000010111","000000000000000000","111111111111111101","111111111111111010","111111111111111111","000000000000000011","000000000000000011","111111111111110100","000000000000001110","000000000000100111","111111111111110110","111111111111010101","111111111111110100","000000000000000010","000000000000010010","000000000000000001","111111111111110101","111111111111110101","000000000000001001","111111111111110001","000000000000000100","111111111111101101","111111111111111010","000000000000010000","000000000000010110","111111111111111011","000000000000000000","111111111111110111","111111111111111101","000000000000011011","111111111111111100","000000000000001011","000000000000101101","111111111111101010","000000000000000100","000000000000100101","000000000000000000","111111111111111111","000000000000001000","000000000000010011","000000000000001010","111111111111101011","111111111111011101","000000000000010000","000000000000001110","000000000000000000","000000000000001011","000000000000001101","111111111111010101","000000000000000111","000000000000101000","000000000000011111","000000000000000111","000000000000010101","111111111111101100","111111111111111010","111111111111110111","111111111111110111","000000000000000011","111111111111111011","000000000000000011","000000000000000000","111111111111101111","111111111111101110","111111111111110100","000000000000010110","000000000000010101","000000000000000000","111111111111111000","000000000000000000","111111111111100101","111111111111101001","000000000000010001","000000000000011011","000000000000000011","111111111111110000","000000000000001111","000000000000000000","111111111111101110","111111111111111101","111111111111010001","000000000000010010","111111111111101001","000000000000011001","111111111111101000","111111111111101101","000000000000001000","000000000000010010","111111111111111000","000000000000010000","111111111111111101","111111111111110010","000000000000000110","000000000000010001","111111111111111010","000000000000001001","000000000000100011","111111111111111101","111111111111110010","000000000000010001","000000000000000000","000000000000001110","000000000000101011","000000000000010001","111111111111101111","111111111111110011","111111111111101100","000000000000001111","000000000000010101","111111111111111101"),
("111111111111111010","000000000000100100","111111111111110100","111111111111100101","111111111110111010","111111111111101100","111111111111110111","111111111111100011","000000000000001100","111111111111110000","000000000000000111","000000000000011100","000000000000110100","111111111111110011","000000000000010010","000000000000000110","111111111111110111","000000000000001000","000000000000010000","000000000000001100","111111111111110000","000000000000010110","000000000000000010","000000000000100101","000000000000010010","111111111111111010","000000000000010000","000000000000001011","111111111111110000","111111111111111011","111111111111111010","000000000000000111","000000000000001111","000000000000000110","000000000000000000","111111111111110001","000000000000000110","000000000000001001","000000000000000110","000000000000011001","000000000000000000","111111111111111111","000000000000000111","111111111111111000","000000000000010001","111111111111100101","111111111111111110","000000000000011110","111111111111111111","111111111111110110","000000000000001010","111111111111101101","000000000000000101","000000000000100001","000000000000010100","000000000000000110","000000000000001001","000000000000000000","000000000000010000","000000000000000001","000000000000000000","111111111111111010","111111111111100111","111111111111111001","111111111111101110","000000000000100001","111111111111100101","000000000000000100","000000000000111110","000000000000000010","111111111111111110","000000000000010100","111111111111011000","111111111111111111","111111111111101100","111111111111111010","000000000000001110","111111111111100000","000000000000000110","000000000000001101","111111111111101110","000000000000010011","000000000000000001","000000000000100011","111111111111110011","111111111111111101","111111111111111110","000000000000000010","111111111111110100","111111111111100011","000000000000100111","111111111111110011","111111111111100001","000000000000000000","111111111111111110","000000000000000110","111111111111000101","000000000000011100","111111111111010111","000000000000010001","111111111111111111","000000000000001110","111111111111111101","111111111111111110","000000000000010001","000000000000010111","111111111111110000","000000000000000000","000000000000010011","000000000000001101","111111111111110011","000000000000010100","000000000000000111","000000000000000001","000000000000100011","111111111111100010","111111111111101101","000000000000010111","000000000000000010","000000000000011111","000000000000001101","000000000000011100","000000000000000010","111111111111101111","111111111111011010","000000000000101010","000000000000101010","111111111111111000"),
("111111111111110110","000000000000011101","000000000000000010","111111111111110011","111111111110101110","111111111111111101","111111111111100111","111111111111111100","111111111111111100","000000000000011101","000000000000010000","000000000000000000","000000000000110000","111111111111110001","000000000000010100","000000000000011000","111111111111110001","000000000000011110","111111111111111111","111111111111111011","000000000000000111","000000000000001100","000000000000000001","000000000000101001","000000000000010000","111111111111111111","111111111111110001","000000000000000110","111111111111111111","111111111111111001","111111111111110111","000000000000000001","000000000000001110","000000000000000000","111111111111111010","000000000000000000","000000000000001011","000000000000001010","000000000000000111","111111111111111000","000000000000100100","000000000000000010","000000000000011110","111111111111110110","111111111111111000","111111111111011111","000000000000000011","111111111111111010","000000000000010001","111111111111110011","000000000000000000","000000000000001001","000000000000010011","000000000000010111","111111111111110001","000000000000001010","111111111111111001","000000000000001100","111111111111111100","111111111111101010","000000000000011001","111111111111011001","000000000000001000","000000000000000010","000000000000000000","000000000000011001","111111111111110001","111111111111111000","000000000000110011","000000000000010000","000000000000001100","000000000000101101","111111111111100000","000000000000010011","000000000000000011","111111111111111010","111111111111101101","111111111111010000","000000000000001110","000000000000000100","000000000000010110","111111111111110000","000000000000001000","111111111111110110","111111111111111100","000000000000001010","111111111111111101","111111111111101100","111111111111111010","111111111111011000","000000000000000110","000000000000001100","111111111111000110","111111111111100100","111111111111110110","000000000000001000","111111111111011100","111111111111111110","000000000000001110","000000000000000010","111111111111110100","111111111111101010","000000000000000000","111111111111111000","000000000000010110","111111111111110010","111111111111110111","000000000000010001","000000000000000100","111111111111101101","000000000000000000","111111111111111010","000000000000000001","111111111111111010","000000000000011000","111111111111111000","000000000000000110","000000000000001101","111111111111111111","000000000000010111","000000000000100011","000000000000001101","000000000000000101","111111111111101001","111111111111011010","000000000000100101","000000000000100001","000000000000000110"),
("000000000000000101","111111111111111100","111111111111111101","111111111111110101","111111111111000010","111111111111111111","111111111111110101","000000000000100010","000000000000010011","000000000000000111","000000000000011101","000000000000000100","000000000000110000","111111111111110010","111111111111101111","000000000000100010","111111111111101110","000000000000011011","111111111111111010","000000000000010101","000000000000010000","111111111111110001","111111111111111001","000000000000001101","000000000000011111","000000000000010001","111111111111010101","000000000000001101","111111111111111011","000000000000000001","111111111111111010","000000000000000110","000000000000000111","111111111111111101","000000000000001010","111111111111110000","111111111111110110","000000000000010010","000000000000010101","111111111111111001","000000000000001000","000000000000000001","000000000000011010","000000000000000001","000000000000000100","111111111111111100","111111111111111110","111111111111010100","111111111111111011","111111111111101110","000000000000011101","111111111111100110","000000000000000010","000000000000101100","000000000000010100","111111111111111001","000000000000000100","111111111111110111","000000000000001100","000000000000001010","000000000000000000","111111111111101100","111111111111100111","000000000000010001","000000000000010110","000000000000000110","000000000000001111","000000000000011010","000000000000011001","000000000000000010","000000000000011110","000000000000101010","111111111111011011","000000000000001010","000000000000010101","111111111111111111","000000000000010011","111111111111110010","111111111111101101","111111111111110001","000000000000001011","000000000000000010","111111111111111010","111111111111111000","000000000000010100","111111111111110001","111111111111101101","111111111111100111","000000000000000100","000000000000010001","000000000000100000","000000000000010000","111111111110111101","000000000000011000","111111111111110001","000000000000001000","111111111111100110","111111111111110110","000000000000000100","000000000000011110","000000000000010111","111111111111011000","111111111111101110","111111111111111000","000000000000010100","000000000000001100","000000000000001110","000000000000010000","111111111111111101","000000000000000000","000000000000010110","111111111111111010","000000000000001010","000000000000001000","000000000000001010","111111111111100011","111111111111110000","000000000000010001","111111111111111001","000000000000011110","000000000000001000","000000000000000100","000000000000000100","111111111111110000","111111111111101111","000000000000001111","000000000000001010","111111111111110111"),
("000000000000011000","111111111111111100","111111111111111110","111111111111101010","000000000000000001","000000000000000100","000000000000001001","000000000000000000","000000000000011101","000000000000000001","000000000000010100","111111111111101100","000000000000010001","111111111111111100","111111111111110111","000000000000110001","111111111111001011","000000000000011101","000000000000000000","000000000000011111","000000000000111000","111111111111110011","111111111111110101","000000000000001111","000000000000010001","000000000000000101","111111111110111001","000000000000011001","111111111111000000","000000000000010001","111111111111111110","111111111111111100","111111111111111001","000000000000010110","000000000000000011","111111111111100110","000000000000000010","000000000000010001","000000000000000011","111111111111101000","000000000000100111","111111111111111111","000000000000010111","000000000000100100","000000000000010010","000000000000010010","000000000000000010","111111111111100100","111111111111110101","111111111111110111","000000000000100011","111111111111101001","111111111111111101","000000000000011100","000000000000100011","000000000000001111","000000000000011011","000000000000000011","000000000000011110","000000000000000010","000000000000011100","111111111111110000","111111111111111011","000000000000000010","000000000000011111","000000000000000000","000000000000100011","111111111111110110","000000000000110010","000000000000000100","000000000000001100","000000000000101101","111111111111111110","000000000000110001","111111111111110001","111111111111111011","111111111111110010","000000000000001011","111111111111111010","000000000000000000","000000000000000110","000000000000001011","111111111111101110","111111111111011010","111111111111110100","000000000000001111","111111111111101101","000000000000000101","000000000000000110","000000000000100011","111111111111111010","000000000000000100","111111111110110100","000000000000010101","000000000000000101","111111111111111010","000000000000010110","000000000000001011","000000000000101011","000000000000001101","111111111111110000","111111111111011100","111111111111111100","000000000000001100","111111111111101100","000000000000001100","000000000000010000","111111111111111011","111111111111011001","000000000000001000","111111111111111001","000000000000011100","000000000000000000","000000000000000001","111111111111111100","111111111111100111","111111111111110001","000000000000011100","111111111111110110","000000000000101001","000000000000101010","111111111111101111","111111111111111110","111111111111101111","111111111111100000","111111111111110110","000000000000011001","000000000000001101"),
("000000000000010000","111111111111101111","000000000000011010","000000000000001011","000000000000110001","111111111111111100","111111111111110110","111111111111111110","000000000000010101","000000000000000001","000000000000001111","111111111111111000","000000000000011011","000000000000000101","111111111111110000","000000000000010101","111111111111011100","000000000000001010","000000000000001100","000000000000011011","000000000000101101","111111111111110011","111111111111111110","000000000000000011","000000000000010111","111111111111101100","111111111111010101","000000000000000110","111111111111011011","000000000000000000","000000000000000001","111111111111111000","000000000000010001","000000000000001010","111111111111110010","000000000000000000","000000000000000111","000000000000000101","111111111111111000","000000000000010010","000000000000011001","000000000000000100","000000000000011101","000000000000100101","000000000000000111","000000000000011101","111111111111100110","111111111111011001","000000000000010011","111111111111110010","000000000000011011","000000000000001101","000000000000000000","000000000000001001","000000000000001000","000000000000001010","000000000000010010","000000000000001110","000000000000001011","000000000000000001","000000000000001000","000000000000011101","000000000000011011","000000000000000000","111111111111111100","111111111111111111","000000000000001010","111111111111110001","000000000000010101","111111111111101100","000000000000001100","000000000000100101","000000000000000010","000000000000100001","111111111111110000","000000000000000101","000000000000000110","000000000000010001","000000000000000101","000000000000000000","000000000000000001","000000000000001111","111111111111100000","000000000000000001","000000000000001000","000000000000000011","111111111111110111","111111111111100110","111111111111110000","000000000000110010","111111111111110101","111111111111111101","111111111110110011","000000000000110100","000000000000011001","000000000000000001","000000000000011100","111111111111110111","000000000000000000","111111111111101101","000000000000001110","000000000000000100","000000000000010110","111111111111101010","111111111111100101","000000000000000010","000000000000010100","000000000000000000","111111111111011010","111111111111111000","111111111111111110","000000000000010011","111111111111100101","000000000000000100","111111111111110101","111111111111110011","111111111111110111","000000000000011110","000000000000000111","000000000000011110","000000000000101110","111111111111100110","111111111111110010","000000000000000001","000000000000000100","000000000000000110","000000000000100011","000000000000001111"),
("000000000000011011","111111111111110011","000000000000010111","111111111111111011","000000000001001001","111111111111110100","000000000000000100","111111111111100110","000000000000010101","111111111111100111","111111111111101001","000000000000010011","000000000000000000","000000000000001001","111111111111101111","000000000000000000","000000000000001100","000000000000011100","000000000000000010","000000000000011011","000000000000110000","111111111111101010","000000000000100000","000000000000000000","000000000000100010","111111111111110001","111111111111011110","000000000000010100","111111111111111000","000000000000010100","000000000000000001","111111111111110011","000000000000010011","111111111111111011","111111111111101111","000000000000001010","000000000000010100","111111111111110101","111111111111111011","000000000000000010","000000000000011011","111111111111010101","000000000000001001","000000000000010011","111111111111111000","000000000000000100","000000000000000000","111111111111111100","000000000000000000","000000000000001110","000000000000001010","111111111111111000","000000000000000111","000000000000001110","000000000000011100","111111111111111110","000000000000001101","000000000000001110","000000000000001101","111111111111110001","000000000000001101","000000000000000010","000000000000100001","111111111111100101","000000000000001000","000000000000000101","000000000000100110","111111111111110000","000000000000010011","111111111111100111","111111111111101111","000000000000001110","000000000000110000","000000000000110100","111111111111110011","111111111111101010","111111111111101100","000000000000001111","000000000000001101","111111111111111010","111111111111101101","000000000000001101","111111111111110011","000000000000010011","111111111111111101","111111111111110011","111111111111111000","111111111111011110","000000000000010100","111111111111111111","111111111111001110","000000000000010101","111111111110111111","000000000000010111","000000000000010101","000000000000001011","000000000000101001","000000000000000110","111111111111110010","111111111111001000","000000000000000010","000000000000000100","000000000000101101","000000000000001011","111111111111111001","111111111111111101","000000000000001100","111111111111110101","000000000000000101","000000000000001111","000000000000000010","000000000000000001","111111111111100111","111111111111110111","000000000000000101","000000000000001111","000000000000010100","111111111111111111","000000000000011010","000000000000100010","000000000000110101","111111111111111001","111111111111101011","000000000000000000","111111111111100001","111111111111110010","000000000000011101","000000000000010011"),
("000000000000001111","111111111111100111","000000000000011111","000000000000100100","000000000000111110","000000000000000001","111111111111101111","111111111111011011","000000000000010010","111111111111100010","000000000000000000","000000000000101001","000000000000000111","000000000000100111","000000000000001011","000000000000010101","000000000000000110","000000000000011010","000000000000010011","000000000000010000","000000000000110000","111111111111100001","000000000000100001","111111111111111010","000000000000100001","000000000000000010","000000000000000110","000000000000010110","000000000000110000","000000000000001011","111111111111110101","111111111111101010","000000000000010101","111111111111101010","111111111111111011","000000000000000000","000000000000011000","111111111111110001","000000000000000000","000000000000001001","000000000000001000","111111111111010010","111111111111111110","000000000000000101","111111111111111000","000000000000000011","111111111111111000","111111111111100111","111111111111111101","000000000000000011","000000000000000011","000000000000001100","000000000000101110","111111111111101111","000000000000010000","111111111111011110","111111111111110110","000000000000100111","000000000000000000","111111111111111000","111111111111111111","000000000000010001","000000000000010011","111111111111111001","000000000000000010","000000000000000001","000000000000101011","111111111111111110","000000000000010101","000000000000000100","000000000000000011","000000000000011110","000000000001000000","000000000000100111","111111111111100001","111111111111110001","111111111111111101","000000000000010100","111111111111110100","000000000000001001","111111111111110100","000000000000000100","111111111111100110","000000000000110000","111111111111111110","000000000000000010","111111111111111110","000000000000000111","111111111111111110","111111111111110100","111111111111011010","000000000000000110","111111111111100001","000000000000000110","000000000000010110","111111111111101110","000000000000011010","111111111111011111","111111111111010001","111111111111001000","000000000000000110","000000000000001000","000000000000011111","000000000000000111","000000000000000000","111111111111111000","000000000000000110","111111111111110101","000000000000001100","000000000000001101","111111111111111101","111111111111111101","111111111111110110","000000000000001010","111111111111101101","000000000000011010","000000000000000101","000000000000000100","000000000000001100","000000000000001001","000000000000010010","111111111111111010","000000000000000000","111111111111111001","111111111111110101","111111111111011110","000000000000011111","000000000000000011"),
("000000000000001000","111111111111110111","000000000000100011","000000000000101011","000000000000011101","111111111111111101","000000000000010100","111111111111111001","000000000000010100","111111111111100001","000000000000001000","000000000000010101","111111111111101011","000000000000100011","111111111111111000","000000000000001010","000000000000001001","000000000000010010","000000000000100111","000000000000100100","000000000000010011","000000000000001110","000000000001000001","000000000000011110","000000000000001110","111111111111101101","000000000000011000","000000000000100100","000000000000100000","111111111111110110","111111111111101101","111111111111110110","000000000000010000","111111111111101001","111111111111111100","000000000000000000","000000000000011001","111111111111111100","000000000000001100","000000000000001001","000000000000011110","111111111111101001","111111111111010001","111111111111100010","111111111111110100","111111111111111111","111111111111101010","111111111111110000","000000000000100010","000000000000100001","000000000000001001","000000000000010010","000000000000001101","111111111111110100","000000000000001101","000000000000000100","111111111111110101","000000000000100001","000000000000001001","000000000000001010","000000000000010111","111111111111111111","000000000000101011","111111111111110011","111111111111111011","000000000000000101","000000000000011010","111111111111110111","000000000000000110","000000000000011101","000000000000001000","000000000000000100","000000000000110010","000000000000100001","111111111111011101","111111111111100110","111111111111100110","000000000000011011","000000000000000110","111111111111110110","000000000000010010","000000000000000000","000000000000000001","000000000000011010","000000000000000011","111111111111110001","111111111111100000","111111111111110110","111111111111101101","111111111111100011","111111111111101111","111111111111111111","111111111111011100","111111111111100111","000000000000110011","111111111111110100","111111111111011111","111111111111111101","111111111111000000","111111111111101111","000000000000000101","000000000000001010","000000000000010010","000000000000001110","000000000000000011","111111111111110110","000000000000010100","111111111111111010","000000000000011101","111111111111110110","000000000000001000","111111111111111100","000000000000000111","000000000000011110","000000000000000110","000000000000100001","111111111111110001","111111111111110101","000000000000000101","000000000000011100","000000000000011011","111111111111111110","111111111111101111","111111111111111001","111111111111101111","111111111111011100","000000000000001011","000000000000011111"),
("000000000000101011","111111111111111001","000000000000001011","000000000000010100","111111111111011101","111111111111111100","000000000000001010","111111111111111110","000000000000001011","111111111111101111","111111111111110111","000000000000011001","000000000000000000","000000000000000000","111111111111111011","000000000000011001","000000000000010100","000000000000011100","000000000000001101","000000000000001111","000000000000010101","111111111111111011","000000000000100111","000000000000010011","000000000000000001","111111111111111011","000000000000001011","000000000000001001","000000000000111000","000000000000011001","111111111111111100","000000000000000100","000000000000000001","111111111111100110","111111111111111011","111111111111111100","000000000000011101","000000000000001010","000000000000001001","000000000000000111","111111111111101101","111111111111000110","111111111111000110","000000000000000011","000000000000000000","111111111111110001","111111111111100011","111111111111101001","000000000000010100","000000000000011001","111111111111101000","000000000000010011","000000000000000110","111111111111110011","000000000000001110","111111111111110111","000000000000010101","000000000000011011","000000000000001001","000000000000010001","000000000000100110","000000000000000000","000000000000110001","111111111111110000","111111111111010001","000000000000001011","000000000000001010","111111111111111011","000000000000001111","000000000000001101","111111111111111110","000000000000011011","000000000000111000","111111111111011110","111111111111101101","111111111111110010","111111111111110101","000000000000001001","000000000000001010","000000000000000000","000000000000010011","111111111111110111","111111111111111010","000000000000010001","000000000000001011","111111111111110111","111111111111101100","000000000000000000","111111111111111100","111111111111100110","111111111111110111","000000000000000000","111111111111010010","000000000000000101","000000000000011110","111111111111101110","111111111111001111","111111111111100010","111111111111001101","000000000000100001","111111111111111000","111111111111111011","000000000000001011","000000000000001000","000000000000010100","000000000000010010","000000000000011000","000000000000001011","000000000000011010","111111111111011010","111111111111111000","000000000000001110","000000000000000010","111111111111111100","111111111111101011","000000000000101111","111111111111101001","111111111111101101","000000000000000011","000000000000010100","000000000000111001","000000000000000111","000000000000000011","000000000000001111","111111111111011101","111111111111100100","000000000000100010","000000000000001010"),
("000000000000011011","000000000000001000","000000000000000010","000000000000011110","111111111111010101","111111111111111000","000000000000000000","000000000000010011","000000000000001001","111111111111101011","000000000000010010","000000000000000110","111111111111110110","000000000000000000","000000000000010011","000000000000000001","111111111111111100","000000000000011000","000000000000101001","000000000000011100","000000000000100111","000000000000011100","000000000000010001","111111111111110000","000000000000010111","111111111111110101","111111111111111101","111111111111111110","000000000000010011","000000000000001011","111111111111110110","111111111111110111","000000000000001100","111111111111011100","000000000000001001","000000000000010110","000000000000010010","000000000000001110","000000000000011100","000000000000010110","000000000000010110","111111111111000111","111111111110110110","111111111111110101","000000000000010011","111111111111101111","000000000000000011","111111111111100101","000000000000000000","000000000000001000","000000000000000000","000000000000010101","000000000000011011","111111111111101110","000000000000000001","000000000000010001","000000000000010100","000000000000010001","111111111111110111","111111111111101100","000000000000011001","000000000000001101","000000000000011110","111111111111110010","111111111111000111","000000000000000010","000000000000010000","000000000000001010","111111111111101111","000000000000000110","000000000000000111","000000000000100110","000000000000001001","111111111110111001","111111111111010010","111111111111111100","111111111111111011","111111111111110101","000000000000000111","000000000000001101","000000000000010100","111111111111110011","000000000000010000","000000000000100100","111111111111110000","111111111111110001","000000000000010000","000000000000001101","111111111111101001","111111111111100010","111111111111110010","000000000000001010","000000000000000011","111111111111101110","111111111111100010","111111111111111111","111111111110111100","111111111111100111","111111111111101001","000000000000101110","111111111111110000","000000000000000101","000000000000010000","000000000000001001","000000000000010101","000000000000001111","000000000000010100","111111111111110000","111111111111110001","111111111111100111","111111111111110110","000000000000010000","111111111111110110","000000000000001011","000000000000010010","000000000000100010","111111111111111111","111111111111111000","000000000000000011","111111111111111111","000000000000110001","000000000000010010","000000000000000011","111111111111110111","111111111111110101","111111111111011001","000000000000010001","000000000000001001"),
("000000000001000111","111111111111111000","000000000000001000","000000000000011110","111111111111001111","000000000000000101","111111111111111010","000000000000010010","111111111111011100","111111111111111110","111111111111110101","000000000000010101","111111111111110011","111111111111110011","000000000000010011","111111111111101100","000000000000000001","000000000000011011","000000000000001111","000000000000000101","000000000000010001","000000000000100101","000000000000011001","111111111111110011","111111111111111111","111111111111111110","000000000000100100","111111111111111111","111111111111001110","000000000000011101","000000000000000110","000000000000001011","000000000000010010","111111111111110011","000000000000001101","000000000000000011","000000000000001110","000000000000001001","000000000000101010","000000000000010100","000000000000000001","111111111111101001","111111111111000111","111111111111101001","000000000000001100","111111111111101100","111111111111101001","111111111111110001","111111111111111000","000000000000001010","000000000000000000","111111111111110101","000000000000011001","111111111111101010","000000000000000101","000000000000000100","000000000000000011","000000000000000100","000000000000010101","000000000000001101","000000000000011010","111111111111100011","000000000000000011","000000000000001110","111111111111011001","000000000000000000","000000000000100001","111111111111111011","111111111111011110","000000000000010000","000000000000001110","000000000000001101","000000000000001111","111111111111000011","111111111111100111","111111111111111101","000000000000000000","000000000000001001","000000000000001100","000000000000010110","000000000000100000","111111111111110010","000000000000001111","000000000000000101","111111111111110100","111111111111111010","111111111111101010","000000000000000001","000000000000001110","111111111110101100","000000000000010011","000000000000000110","111111111111111011","111111111111111001","111111111111100011","111111111111111011","111111111111000101","111111111111111100","111111111111111110","000000000000101101","000000000000000000","111111111111111111","000000000000000111","000000000000001001","111111111111111111","111111111111110000","111111111111111110","111111111111111110","111111111111101111","111111111111111000","000000000000001001","000000000000000001","111111111111101111","111111111111110101","000000000000011000","000000000000000111","111111111111110000","111111111111111111","111111111111110110","111111111111110001","000000000000011011","000000000000010100","111111111111101001","000000000000000010","111111111111100000","111111111111111000","000000000000001000","111111111111111000"),
("000000000000011101","111111111111101100","111111111111111010","000000000000010111","111111111111000111","111111111111111110","111111111111111000","000000000000010111","111111111111110101","111111111111110101","000000000000001100","000000000000000000","111111111111101111","000000000000001000","111111111111101110","000000000000001010","000000000000001001","000000000000101001","000000000000110110","000000000000100010","000000000000100011","000000000000011000","000000000000011000","111111111111111000","000000000000000000","000000000000001010","000000000000101000","111111111111101110","111111111111000101","000000000000001100","111111111111101110","111111111111101010","000000000000001111","111111111111101011","000000000000010000","111111111111111001","000000000000010100","000000000000000001","000000000000101001","000000000000001010","000000000000000010","111111111111010111","111111111111010011","111111111111011001","000000000000000010","111111111111010110","111111111111100100","111111111111100101","000000000000011110","000000000000000100","111111111111111000","000000000000100001","111111111111101111","111111111111101010","000000000000000110","000000000000010110","000000000000001101","000000000000010000","000000000000010101","111111111111101110","000000000000100110","000000000000010000","111111111111100011","111111111111111111","000000000000000101","111111111111101000","000000000000011010","111111111111101101","111111111111110011","000000000000011101","000000000000001000","000000000000101000","000000000000101001","111111111110110100","111111111111101001","111111111111101011","111111111111111100","000000000000000000","111111111111111010","000000000000001100","111111111111110010","111111111111111110","111111111111101001","111111111111111101","000000000000001110","000000000000000001","111111111111111010","111111111111101101","111111111111110010","111111111111011111","111111111111111110","000000000000010111","111111111111110001","000000000000000011","111111111111101010","111111111111111110","111111111111011110","000000000000000010","000000000000000011","000000000000101001","111111111111101100","111111111111110000","000000000000010110","111111111111111001","000000000000000010","111111111111111010","111111111111111101","000000000000001001","111111111111110101","111111111111101110","111111111111110111","111111111111101000","000000000000001011","111111111111110111","000000000000110101","000000000000101010","000000000000001010","000000000000000000","111111111111111100","000000000000010101","000000000000010010","111111111111110101","111111111111110000","000000000000010110","000000000000000000","111111111111001110","000000000000011010","000000000000001101"),
("000000000000101100","111111111111111001","111111111111110110","111111111111110101","111111111111100011","111111111111111010","000000000000000000","111111111111110111","111111111111111111","000000000000000000","000000000000100010","111111111111111110","111111111111110001","111111111111110011","111111111111101100","000000000000001100","111111111111101100","000000000000011100","000000000000001101","000000000000000001","000000000000011111","000000000000010100","000000000000000111","000000000000010010","000000000000001001","000000000000000001","000000000000001010","111111111111100000","111111111111000101","000000000000000100","111111111111101111","111111111111100011","000000000000011010","111111111111100111","000000000000001110","111111111111101000","000000000000100000","000000000000001100","000000000000001011","000000000000011111","000000000000000011","111111111111101111","111111111111000010","111111111111010010","111111111111111101","111111111111101110","111111111111100110","111111111111100110","000000000000101010","111111111111101101","000000000000101101","000000000000101011","000000000000100001","111111111111011000","111111111111100100","000000000000000011","000000000000010100","111111111111110001","000000000000011000","000000000000010001","000000000000010010","000000000000001110","111111111111010100","000000000000000011","111111111111101110","000000000000000000","000000000000011100","111111111111101110","111111111111101001","000000000000011100","000000000000000000","000000000000011111","000000000000101000","111111111111001111","111111111111000010","111111111111011110","000000000000011001","111111111111111110","000000000000000011","000000000000010111","111111111111110000","000000000000001010","000000000000000100","000000000000000000","111111111111111101","111111111111100101","000000000000001010","111111111111111011","111111111111100101","111111111111101010","000000000000011100","111111111111101101","111111111111110110","111111111111111111","111111111111110101","111111111111100110","111111111111011111","111111111111110111","111111111111110100","000000000000010001","000000000000000000","000000000000000000","111111111111110011","000000000000011000","000000000000101001","000000000000001000","111111111111011110","111111111111111000","111111111111101011","111111111111110000","000000000000000111","111111111111101111","111111111111111111","000000000000001001","000000000000011001","000000000000000100","111111111111101000","000000000000001010","111111111111111010","111111111111100101","000000000000011001","000000000000001011","111111111111100101","000000000000010010","111111111111110001","111111111111100110","000000000000100001","111111111111101110"),
("000000000001000101","000000000000011101","000000000000100110","111111111111101011","111111111111010100","111111111111101111","111111111111110111","111111111111111110","111111111111011010","000000000000000001","111111111111101101","000000000000001010","111111111111011110","111111111111101010","111111111111100100","000000000000000000","111111111111000101","000000000000001110","000000000000000000","111111111111011110","000000000000011101","000000000000001101","111111111111101100","000000000000011100","000000000000011000","111111111111100100","000000000000100101","111111111111001000","111111111111010010","000000000000000010","000000000000011110","111111111111001010","111111111111111010","111111111111111011","000000000000001000","111111111111010010","000000000000100100","000000000000011001","000000000000101001","000000000000001111","000000000000000101","111111111111111101","111111111111100101","111111111111101000","000000000000001101","111111111111111000","111111111111100101","111111111111110000","000000000000101010","111111111111011010","000000000000001000","000000000000101001","000000000000000101","111111111111111001","111111111111111011","000000000000010110","000000000000101011","111111111111101110","111111111111101101","111111111111111110","000000000000011110","111111111111100111","111111111110100001","111111111111111001","000000000000001000","000000000001000101","000000000000011010","111111111111011101","111111111111110011","000000000000100011","111111111111100101","111111111111110011","000000000000110100","111111111111010110","111111111110110000","111111111111111010","000000000000010001","111111111111011100","000000000000001000","111111111111100110","000000000000010010","000000000000011001","111111111111101111","111111111111001101","111111111111111101","111111111111100000","000000000000010000","000000000000000011","111111111111111010","111111111111101101","000000000000011111","000000000000011101","000000000000010110","111111111111011100","111111111111100011","111111111111010000","111111111111011010","111111111111100010","000000000000010110","111111111111111111","111111111111111001","000000000000001101","111111111111110011","000000000000011010","000000000000011000","111111111111111001","000000000000011011","111111111111110001","000000000000000101","111111111111111010","000000000000100000","111111111111101010","000000000000000000","111111111111101001","000000000000110011","111111111111011000","111111111111101100","000000000000001110","000000000000010101","000000000000000001","111111111111110111","000000000000100100","111111111111011111","111111111111110001","111111111111011100","111111111111100100","000000000000000111","000000000000010111"),
("000000000000110001","000000000000011100","000000000000110111","111111111111111000","111111111111011100","111111111111111000","000000000000000001","111111111111111011","000000000000001100","111111111111110110","111111111111100001","000000000000010001","111111111111101100","111111111111101001","111111111111100000","111111111111010010","111111111111011011","111111111111110000","111111111111101010","111111111111110011","000000000000000000","111111111111011100","111111111111010101","000000000000001001","000000000000100000","111111111111101100","000000000000100011","111111111111001000","111111111111010101","000000000000100000","000000000000101100","111111111110111000","111111111111110100","000000000000000011","000000000000011100","000000000000010111","000000000000000111","000000000000110010","000000000000011100","000000000000100111","000000000000011101","000000000000001000","111111111111110011","111111111111110010","000000000001010000","111111111111101110","000000000000001010","000000000000101101","000000000000011111","111111111111001100","111111111111110011","000000000000101100","111111111111101000","000000000000001100","000000000000000000","000000000000011111","000000000000100000","111111111111010101","111111111111011100","000000000000001011","111111111111111010","111111111111011100","111111111111000111","111111111111111011","000000000000000101","000000000000110110","000000000000010000","000000000000000100","111111111111011101","000000000000001010","111111111111100010","111111111111111011","000000000000010000","111111111111101001","111111111111110001","000000000000001000","000000000000101110","111111111111100110","111111111111110011","111111111111111101","000000000000010110","000000000001001010","000000000000001000","111111111111001101","111111111111110101","111111111111111110","000000000000001100","000000000000011110","111111111111111101","111111111111011000","000000000000001100","111111111111101010","111111111111111010","111111111111010010","111111111111101100","111111111111101101","000000000000001001","111111111111111100","000000000000001101","000000000000011110","000000000000111010","000000000000001010","111111111111011100","000000000000000110","000000000000010011","000000000000000100","000000000000000010","000000000000000000","000000000000010011","111111111111110001","000000000000100100","000000000000001100","000000000000010001","000000000000001110","000000000000010010","111111111111000010","111111111111100111","111111111111110110","000000000000101101","111111111111111111","000000000000001010","000000000000101010","111111111111100101","111111111111011010","111111111111011110","111111111111101100","000000000000010010","000000000000110001"),
("111111111111111000","111111111111110100","000000000000001010","000000000000000000","111111111111110111","000000000000010101","000000000000000111","111111111111110000","000000000000011000","111111111111011101","111111111111111110","000000000000010000","000000000000011011","111111111111011000","000000000000000000","000000000000001101","111111111111010001","000000000000000101","000000000000001011","111111111111111111","111111111111111111","111111111111110100","111111111111000100","000000000000001100","000000000000000000","000000000000100001","000000000000101010","111111111111100011","111111111111110000","000000000000001010","111111111111111111","111111111111110011","111111111111110010","000000000000001001","000000000000101000","000000000000011000","111111111111110101","000000000000100001","000000000000011011","000000000000000010","000000000000001011","000000000000011000","111111111111111111","111111111111111111","000000000000111010","000000000000001101","000000000000010000","111111111111111111","000000000000101000","111111111111101110","111111111111110101","000000000000010110","111111111111101111","111111111111111101","000000000000001011","000000000000010100","000000000000100101","111111111111110101","000000000000000110","111111111111111111","000000000000000011","000000000000001010","111111111111101110","000000000000010101","111111111111000000","111111111111111010","000000000000000110","111111111111110111","111111111111111011","000000000000100100","000000000000000010","000000000000011110","111111111111110110","111111111111110001","000000000000000101","000000000000001000","000000000000101101","000000000000000111","111111111111111100","000000000000001000","000000000000001010","000000000000011100","111111111111110110","111111111111011011","000000000000010101","111111111111011100","000000000000000001","000000000000101001","000000000000001011","111111111111100011","000000000000000011","111111111111110100","000000000000000111","111111111111010010","000000000000011101","000000000000001010","000000000000000010","111111111111101001","111111111111101010","000000000000011001","000000000000011010","000000000000011011","111111111111110100","000000000000100001","000000000000100100","000000000000010100","000000000000100011","000000000000010010","111111111111111000","111111111111101100","000000000000011101","000000000000001001","000000000000011010","111111111111111111","000000000000011111","111111111111101000","111111111111100110","111111111111111000","000000000000110111","000000000000011010","000000000000001011","000000000000000010","111111111111011100","111111111111011000","111111111111100010","000000000000001010","000000000000000111","000000000000001000"),
("000000000000001100","111111111111111110","000000000000000001","000000000000000100","111111111111111000","111111111111100101","000000000000001111","111111111111111110","000000000000001010","111111111111111010","000000000000100001","000000000000011110","000000000000000110","111111111111110001","111111111111111000","111111111111110101","000000000000000011","000000000000010001","000000000000011001","000000000000000000","000000000000110000","000000000000010100","111111111111111101","000000000000000110","000000000000100110","000000000000000000","000000000000001001","111111111111011010","111111111111111100","111111111111111111","000000000000101001","000000000000000111","000000000000000000","000000000000001001","000000000000101100","000000000000000101","000000000000000000","111111111111111111","111111111111110110","111111111111101011","000000000000010111","000000000000101110","111111111111100100","111111111111100110","000000000000001010","000000000000000110","000000000000010100","000000000000100101","000000000000011111","111111111111111010","000000000000010011","000000000000100010","000000000000010101","111111111111111111","000000000000001100","000000000000001100","000000000000001010","111111111111110000","000000000000010000","000000000000000011","000000000000000111","000000000000000100","111111111111101100","111111111111111001","111111111111111000","000000000000010011","000000000000010101","000000000000100001","000000000000000001","000000000000001010","000000000000000000","000000000000100100","000000000000010000","000000000000000110","111111111111101101","111111111111111000","000000000000001000","111111111111101001","111111111111101110","000000000000000011","111111111111111011","000000000000010100","000000000000000100","111111111111101110","000000000000001000","111111111111101010","111111111111111111","000000000000001001","111111111111110000","111111111111110111","111111111111101111","000000000000100010","000000000000011000","111111111111001111","000000000000000110","111111111111111011","111111111111110100","000000000000000001","111111111111111011","111111111111111010","111111111111111111","000000000000100010","111111111111111110","000000000000100110","000000000000101000","000000000000010010","000000000000000101","000000000000010010","111111111111010101","111111111111101101","000000000000011010","000000000000001001","000000000000010110","000000000000000000","000000000000001011","111111111111110100","000000000000000011","000000000000011001","000000000000011110","000000000000000110","000000000000000101","000000000000000101","111111111111110000","111111111111110001","111111111111111101","111111111111111011","000000000000100001","000000000000001100"),
("000000000000001000","111111111111110100","000000000000000110","000000000000001000","000000000000000110","111111111111100011","000000000000001100","111111111111101010","111111111111111011","000000000000011001","000000000000000000","111111111111110100","111111111111111010","000000000000001110","000000000000000111","111111111111111101","111111111111101011","111111111111110101","000000000000011010","000000000000010100","000000000000011100","111111111111110110","111111111111110101","000000000000000111","000000000000001001","000000000000001001","111111111111111101","000000000000010000","111111111111111001","000000000000001001","000000000000000000","111111111111111111","000000000000001110","111111111111110111","000000000000011010","111111111111101001","000000000000011100","111111111111101000","111111111111110010","000000000000000110","000000000000000000","111111111111111110","111111111111111001","000000000000000000","111111111111100110","000000000000000101","111111111111110110","111111111111111011","000000000000001000","000000000000010110","111111111111111100","000000000000001001","000000000000001101","000000000000001011","000000000000010010","000000000000001001","111111111111110111","000000000000001100","000000000000001000","000000000000000001","000000000000000000","000000000000000101","111111111111110111","111111111111100111","000000000000000011","000000000000001010","111111111111111100","111111111111111111","111111111111111111","000000000000001000","111111111111111111","111111111111111111","000000000000000110","000000000000011001","111111111111110111","000000000000000000","000000000000001001","000000000000001100","000000000000100000","111111111111111010","000000000000000111","111111111111101011","111111111111110101","000000000000001110","111111111111110101","111111111111111000","111111111111111011","111111111111110001","000000000000000101","000000000000010000","111111111111110111","111111111111101101","000000000000000111","111111111111110100","000000000000010101","000000000000001000","111111111111100100","000000000000000000","111111111111111111","000000000000001111","111111111111110010","111111111111111010","111111111111111000","111111111111100100","000000000000010010","111111111111110001","111111111111110101","000000000000001001","111111111111101000","000000000000000101","000000000000011001","111111111111111010","111111111111101001","000000000000001110","000000000000001001","000000000000000110","111111111111110000","000000000000001111","111111111111111000","000000000000010000","000000000000010011","111111111111111011","111111111111110011","000000000000011000","000000000000010101","111111111111111110","000000000000000000","000000000000000000"),
("111111111111111111","000000000000000001","000000000000010111","000000000000001010","000000000000010110","000000000000000001","111111111111111000","111111111111011110","000000000000011101","000000000000011111","111111111111110111","111111111111111111","000000000000000110","000000000000011100","000000000000010100","000000000000000001","000000000000001000","000000000000010011","000000000000001110","000000000000011011","000000000000001010","000000000000010010","000000000000001010","111111111111101000","000000000000010001","000000000000000100","000000000000010001","000000000000000000","000000000000010101","000000000000100011","111111111111100001","111111111111111111","111111111111101000","000000000000000011","000000000000010011","111111111111011000","000000000000011010","000000000000000000","111111111111111100","000000000000000011","111111111111111010","000000000000100110","000000000000100000","000000000000000100","111111111111101111","000000000000001101","000000000000001110","000000000000000101","000000000000010110","000000000000010000","111111111111110011","111111111111101100","000000000000011110","000000000000000111","000000000000000001","000000000000001011","111111111111111011","000000000000001000","000000000000001000","000000000000001101","000000000000011111","000000000000010000","111111111111110101","111111111111111011","111111111111010100","000000000000010110","111111111111101101","111111111111101010","111111111111110011","000000000000101011","111111111111101011","000000000000010111","111111111111101111","000000000000010001","111111111111100010","000000000000001001","111111111111111100","000000000000000010","111111111111111010","000000000000000101","111111111111101011","111111111111110000","111111111111100111","000000000000100100","111111111111110111","000000000000101000","000000000000001110","111111111111111111","111111111111111110","111111111111111010","000000000000010001","000000000000000101","000000000000100001","111111111111101010","000000000000001101","000000000000001000","000000000000000010","111111111111101100","000000000000001011","000000000000001101","111111111111100010","111111111111101000","111111111111111101","111111111111111011","111111111111111011","111111111111100111","111111111111110100","000000000000000000","111111111111110001","000000000000010110","000000000000000110","111111111111101001","111111111111110000","111111111111111100","000000000000000110","111111111111011100","111111111111101000","000000000000010100","111111111111101001","000000000000000001","000000000000010010","111111111111101110","000000000000101000","000000000000101011","000000000000011000","111111111111011101","000000000000010110","000000000000000101"),
("000000000000001100","000000000000001001","000000000000000101","111111111111100101","000000000000000101","111111111111101111","111111111111110110","111111111111101100","111111111111101111","000000000000000000","000000000000000100","111111111111111100","111111111111101000","000000000000000001","000000000000010100","111111111111100100","000000000000001011","111111111111100101","000000000000010110","000000000000001111","111111111111101010","000000000000010110","000000000000100000","000000000000001010","111111111111111101","111111111111101110","000000000000011101","111111111111101100","000000000000001110","111111111111110010","111111111111100110","000000000000001011","000000000000001010","111111111111101100","111111111111111011","000000000000011001","111111111111111000","000000000000001101","000000000000000111","000000000000001001","111111111111101011","111111111111111110","000000000000010000","111111111111111000","111111111111111010","111111111111110010","000000000000001000","000000000000000101","000000000000001111","000000000000100010","111111111111111011","000000000000000010","000000000000001100","111111111111110010","000000000000000001","000000000000000101","000000000000000010","000000000000010100","111111111111111100","000000000000000101","111111111111111100","111111111111111000","111111111111101111","111111111111111001","111111111111001010","111111111111110000","111111111111111000","111111111111110100","000000000000011101","111111111111101111","111111111111110001","000000000000001011","111111111111011010","111111111111101111","111111111111111000","111111111111110001","000000000000001101","111111111111110101","000000000000001110","000000000000101100","111111111111101110","111111111111101111","111111111111101001","000000000000010011","000000000000001101","000000000000010110","111111111111110101","111111111111110100","000000000000001001","000000000000000101","111111111111101010","111111111111110110","111111111111110111","111111111111110011","111111111111110011","000000000000000000","000000000000000010","111111111111101111","111111111111111011","111111111111100010","000000000000001100","111111111111111010","000000000000011000","111111111111111110","000000000000011101","000000000000000000","000000000000000000","000000000000000110","000000000000101001","111111111111110101","000000000000000100","111111111111110000","111111111111111001","000000000000010010","000000000000100011","111111111111101001","111111111111101111","000000000000001001","000000000000000001","111111111111110000","000000000000000101","000000000000001110","111111111111101110","111111111111110001","111111111111111101","111111111111011111","111111111111100101","111111111111111000"),
("000000000000000101","000000000000000101","111111111111101111","000000000000000110","000000000000001010","111111111111100100","111111111111110001","111111111111011011","000000000000101010","000000000000000010","000000000000011000","111111111111110001","000000000000000100","000000000000000101","111111111111110101","111111111111111110","000000000000001001","000000000000000010","000000000000001000","000000000000011011","000000000000010001","000000000000010010","000000000000001101","111111111111111101","000000000000000011","000000000000001100","000000000000001111","000000000000001100","000000000000100011","111111111111100011","111111111111011001","000000000000000100","000000000000000001","000000000000000001","000000000000010110","000000000000001000","111111111111111101","111111111111110100","111111111111101111","111111111111110111","111111111111111011","111111111111111000","000000000000011111","000000000000011101","111111111111110111","000000000000000111","000000000000011110","111111111111011011","000000000000011000","000000000000000000","000000000000101100","000000000000000101","000000000000001101","111111111111101010","000000000000000000","000000000000010110","111111111111100000","000000000000011001","111111111111111110","000000000000000001","111111111111111011","111111111111111010","111111111111010110","000000000000001001","111111111111100111","000000000000000011","000000000000001100","000000000000000010","000000000000000011","111111111111100010","000000000000010000","000000000000000100","111111111111101000","000000000000011100","111111111111110011","111111111111110111","000000000000000000","000000000000011001","000000000000000110","000000000000010000","111111111111100111","000000000000000001","000000000000000000","000000000000010011","000000000000010010","000000000000010001","111111111111111011","111111111111111101","111111111111111100","000000000000010110","111111111111001110","111111111111011010","111111111111110111","000000000000011101","000000000000001100","111111111111101100","000000000000011111","111111111111101101","000000000000011010","111111111111110100","111111111111110111","111111111111101111","111111111111111010","000000000000000101","000000000000010001","000000000000011100","111111111111110001","111111111111110001","000000000000011001","000000000000001010","111111111111110101","000000000000001001","000000000000010000","000000000000010101","000000000000010010","000000000000001111","000000000000011011","000000000000011000","111111111111101111","000000000000001011","000000000000010010","000000000000000001","000000000000010011","111111111111111001","000000000000001001","111111111111010010","000000000000000000","000000000000000101"),
("111111111111100010","000000000000011010","000000000000010010","111111111111111101","000000000000000111","111111111111110011","111111111111110000","000000000000001110","000000000000000011","000000000000011111","000000000000001100","000000000000001001","000000000000001100","000000000000001110","000000000000000010","111111111111110101","000000000000000000","111111111111101110","000000000000000110","000000000000000100","111111111111111100","000000000000101001","000000000000100010","111111111111100000","111111111111110111","000000000000000000","000000000000010111","000000000000000010","000000000000010001","000000000000000000","111111111111100010","000000000000100100","111111111111011110","111111111111111100","111111111111100000","111111111111111001","111111111111110001","000000000000010110","000000000000010000","111111111111111110","000000000000000100","111111111111010100","000000000000011100","000000000000010010","111111111111111111","000000000000010101","000000000000100111","111111111110101110","000000000000000001","000000000000001010","000000000000000011","111111111111111111","000000000000000011","111111111111111011","111111111111111010","111111111111111001","111111111111010111","000000000000001011","000000000000001001","000000000000001101","111111111111100010","111111111111110011","111111111111011100","111111111111101110","000000000000001000","000000000000000100","111111111111100100","111111111111100101","000000000000010011","111111111111111001","000000000000001001","000000000000010110","000000000000001000","000000000000100111","000000000000001110","000000000000000011","000000000000000000","111111111111110001","000000000000001111","111111111111111010","111111111111100100","111111111111100110","111111111111011011","111111111111110001","111111111111111111","000000000000010001","000000000000011110","000000000000010101","111111111111101011","000000000000100001","111111111111100101","111111111111010110","000000000000001110","111111111111101110","111111111111110011","111111111111101111","000000000000001011","000000000000000000","000000000000010001","111111111111011000","000000000000000001","111111111111101001","111111111111111100","111111111111101011","000000000000011000","111111111111111101","111111111111110100","000000000000101000","000000000000011001","111111111111101011","111111111111101011","000000000000001100","111111111111111010","000000000000000000","000000000000001100","000000000000010011","000000000000000111","000000000000101010","111111111111001110","111111111111111110","000000000000001111","111111111111101101","111111111111101010","000000000000010001","000000000000000111","111111111111010001","111111111111111111","111111111111110101"),
("111111111111001110","000000000000010101","000000000000010001","111111111111101011","000000000000011011","111111111111100111","000000000000001001","000000000000111011","000000000000010101","111111111111101110","000000000000001010","111111111111111010","000000000000010110","111111111111111010","000000000000001101","000000000000000011","111111111111101110","111111111111111000","000000000000001010","111111111111110111","111111111111110000","000000000000001000","111111111111110110","111111111111100001","000000000000001010","111111111111110000","000000000000001001","111111111111111010","000000000000000110","111111111111101000","111111111111110101","111111111111110000","111111111111111111","111111111111010010","111111111111100100","000000000000010011","000000000000010010","000000000000011100","000000000000000000","000000000000001111","000000000000001100","111111111111010110","000000000000010111","111111111111111000","000000000000010010","111111111111110001","000000000000010110","111111111111100011","000000000000000000","000000000000000111","111111111111111100","111111111111100111","111111111111111101","000000000000011001","000000000000010001","000000000000011100","111111111110111100","111111111111110100","111111111111110110","111111111111101101","000000000000000110","111111111111011000","111111111111101101","111111111111101001","111111111110111101","111111111111111110","111111111111101100","111111111111100011","000000000000001000","111111111111101010","111111111111110001","111111111111110000","000000000000011100","000000000000000010","111111111111110110","000000000000010010","111111111111111011","111111111111101011","000000000000100000","111111111111110100","111111111111100000","000000000000001110","111111111111010010","111111111111011001","111111111111110101","000000000000001011","111111111111110101","111111111111101011","111111111111011001","111111111111111100","111111111111010100","111111111111100110","000000000000010110","111111111111101111","000000000000001101","111111111111110110","111111111111100000","000000000000100001","111111111111001110","000000000000000001","111111111111100000","111111111111011101","111111111111111000","000000000000000010","000000000000001111","000000000000001011","000000000000010010","000000000000011000","111111111111100110","000000000000000101","000000000000000110","000000000000001101","000000000000001101","111111111111111011","000000000000010010","111111111111110011","111111111111111001","000000000000100001","111111111111100110","000000000000000001","000000000000010101","111111111111110100","111111111111111011","000000000000100110","000000000000001001","111111111111011001","111111111111111010","111111111111101100"),
("111111111111000100","000000000000100001","111111111111111110","111111111111100111","111111111111111001","111111111111011100","000000000000011011","111111111111111110","000000000000001011","111111111111010000","000000000000000000","000000000000001001","000000000000001110","000000000000001000","000000000000000011","111111111111011110","111111111111010011","000000000000000100","000000000000000111","000000000000001011","111111111111111110","000000000000001011","111111111111110000","111111111111100111","111111111111110110","111111111111111000","000000000000000001","111111111111110001","111111111111110010","111111111111101110","000000000000000000","111111111111111000","000000000000010000","111111111111110100","111111111111110001","000000000000001001","000000000000010011","000000000000011001","111111111111110010","000000000000001110","000000000000001010","111111111111110111","111111111111110010","000000000000000010","000000000000001000","000000000000001000","000000000000001000","111111111111101111","000000000000010100","000000000000001011","111111111111110001","111111111111101111","000000000000000000","000000000000101011","111111111111110100","000000000000010001","111111111111011100","000000000000011001","000000000000011110","111111111111110001","111111111111101101","111111111111010010","111111111111101101","111111111111101111","111111111111000010","000000000000001110","111111111111011010","111111111111111011","000000000000011101","111111111111101011","000000000000010001","000000000000001101","111111111111110101","000000000000001001","000000000000011000","000000000000001001","000000000000000001","111111111111100110","000000000000010100","000000000000001010","000000000000001001","111111111111111101","111111111111011100","111111111111011011","111111111111110101","111111111111100000","111111111111111110","111111111111111101","111111111111110001","000000000000000101","111111111111011101","111111111111111000","000000000000010110","111111111111111110","000000000000011110","111111111111101101","111111111111100111","000000000000000000","111111111111101111","000000000000010101","111111111111011001","000000000000011100","111111111111010101","000000000000000010","111111111111110111","000000000000010001","000000000000010000","000000000000001111","000000000000011000","111111111111100110","000000000000001100","000000000000010110","111111111111110101","000000000000010000","000000000000010011","111111111111010100","111111111111111110","111111111111111111","111111111111101010","111111111111111001","000000000000000100","111111111111110100","111111111111111100","000000000000000011","111111111111101011","111111111111111101","111111111111110101","000000000000010001"),
("111111111110110001","000000000000001100","000000000000000111","000000000000000010","000000000000010010","111111111111111101","111111111111110011","111111111111110001","111111111111111101","111111111111111110","000000000000100011","000000000000101100","000000000000011010","000000000000010101","000000000000000111","111111111111111110","111111111111100000","000000000000001001","111111111111111110","111111111111110110","000000000000000111","000000000000010001","111111111111111011","111111111111110111","111111111111110101","000000000000001010","000000000000001000","000000000000000001","111111111111110000","111111111111010010","111111111111101011","000000000000000110","111111111111110100","111111111111101010","000000000000001011","000000000000010000","111111111111111101","000000000000001011","111111111111110001","111111111111111011","000000000000011011","111111111111100111","000000000000011110","111111111111101001","000000000000000000","111111111111111110","000000000000001110","000000000000001001","000000000000001100","000000000000010001","111111111111111110","111111111111110010","111111111111111111","000000000000011000","000000000000001100","000000000000000001","111111111111100000","000000000000000011","000000000000010111","111111111111110111","111111111111110000","111111111111010010","111111111111101011","000000000000000100","111111111111011000","000000000000011100","111111111111011101","000000000000010100","000000000000110000","000000000000000010","111111111111111111","000000000000001111","111111111111010111","000000000000001101","000000000000001111","000000000000010010","111111111111100000","111111111111110101","000000000000001000","111111111111011110","000000000000001010","000000000000000001","111111111111101110","000000000000001000","000000000000001110","000000000000000000","000000000000010010","111111111111110111","111111111111110011","000000000000000111","111111111111011011","000000000000001100","000000000000001100","111111111111110111","000000000000010100","111111111111111000","111111111111100110","111111111111101111","111111111111111011","000000000000000001","111111111111110100","000000000000000111","111111111111011110","111111111111111100","111111111111100001","111111111111111000","000000000000011000","000000000000001101","000000000000001000","000000000000000010","000000000000001010","000000000000000011","000000000000010011","000000000000010101","000000000000011010","111111111111111100","111111111111110001","000000000000000000","111111111111101001","000000000000100010","111111111111111011","111111111111100111","000000000000000001","000000000000001111","111111111111111010","000000000000010011","000000000000010001","111111111111111101"),
("111111111111010101","000000000000000000","000000000000000111","111111111111101010","000000000000110111","111111111111111011","000000000000000100","000000000000011010","000000000000000110","111111111111101101","000000000000100101","000000000000001111","000000000000010011","000000000000010111","000000000000010100","000000000000000100","111111111111011000","111111111111111101","000000000000010101","111111111111111101","111111111111101011","000000000000010011","000000000000000010","111111111111011001","111111111111111011","000000000000000110","000000000000010100","000000000000011100","111111111111011100","111111111111110110","000000000000001101","000000000000000000","111111111111101111","111111111111110111","000000000000000100","000000000000000000","111111111111110100","111111111111110111","000000000000010001","000000000000001011","000000000000010100","111111111111110010","000000000000000110","000000000000000000","000000000000001000","111111111111110001","111111111111111111","111111111111110001","000000000000001000","000000000000010010","111111111111100101","111111111111110011","111111111111110100","000000000000100011","000000000000000011","111111111111110111","000000000000001011","000000000000001101","000000000000011000","111111111111110110","111111111111101100","111111111111011100","111111111111101011","111111111111101111","111111111111110110","000000000000000111","111111111111011101","111111111111110100","000000000000101110","000000000000000010","111111111111110101","000000000000011001","111111111111011111","111111111111101111","111111111111111110","000000000000011010","111111111111111100","000000000000000011","000000000000000100","111111111111110010","111111111111110110","111111111111111101","111111111111010110","111111111111111110","000000000000011010","111111111111101111","000000000000011000","111111111111110001","000000000000000011","111111111111010000","111111111111100011","000000000000010101","000000000000001011","000000000000000000","000000000000000011","111111111111101001","111111111111101011","000000000000001001","111111111111100111","000000000000011011","111111111111100010","000000000000100110","111111111111100101","111111111111111000","111111111111110010","000000000000001011","000000000000010100","000000000000011100","000000000000000000","111111111111111100","000000000000010100","111111111111111110","000000000000001110","000000000000000110","000000000000001101","111111111111111011","000000000000001011","000000000000011110","000000000000000000","000000000000100110","000000000000000110","111111111111110100","000000000000001000","000000000000000001","111111111111110011","000000000000001110","000000000000011000","000000000000000010"),
("111111111111100111","000000000000000111","000000000000001000","111111111111101100","000000000000100000","111111111111110000","111111111111111011","000000000000011010","000000000000000110","111111111111101111","000000000000011101","000000000000100100","000000000000101000","000000000000001101","000000000000001111","000000000000001110","111111111111011001","000000000000001111","111111111111111001","111111111111011111","111111111111110010","000000000000000011","000000000000010001","111111111111010101","111111111111110110","111111111111111000","000000000000010000","000000000000001010","111111111111110100","111111111111011000","111111111111111010","111111111111111111","111111111111110100","000000000000001111","000000000000011000","111111111111111111","111111111111111100","111111111111011110","111111111111111111","000000000000000100","000000000000001101","111111111111110101","000000000000100101","000000000000001100","111111111111101101","111111111111101010","000000000000001000","000000000000000001","111111111111111001","111111111111111101","111111111111110000","000000000000000010","000000000000001001","000000000000101000","111111111111101111","000000000000010110","000000000000000000","000000000000000100","000000000000010001","111111111111111110","000000000000000011","111111111111010100","111111111111110100","000000000000010001","111111111111111010","000000000000010011","111111111111100011","000000000000000101","000000000001001001","111111111111111010","111111111111111111","111111111111111001","111111111111101011","000000000000000010","111111111111101000","111111111111110000","000000000000001000","111111111111101101","000000000000001111","000000000000000010","111111111111111000","000000000000000000","111111111111111101","000000000000101110","000000000000000111","111111111111101100","000000000000001010","111111111111111100","111111111111111010","111111111111000011","000000000000000000","000000000000010101","000000000000100100","111111111111111010","111111111111111111","000000000000011000","111111111111000011","000000000000010011","111111111111011001","000000000000001100","111111111111101111","000000000000101011","111111111111110001","000000000000010000","000000000000000001","111111111111111001","000000000000010001","000000000000010000","000000000000001010","000000000000000000","000000000000000000","000000000000100010","111111111111110000","000000000000000110","000000000000001001","000000000000000100","000000000000000111","000000000000001101","000000000000001110","111111111111111111","111111111111111011","111111111111111110","111111111111111111","111111111111111010","111111111111100110","000000000000001100","000000000000010100","000000000000001010"),
("000000000000010100","000000000000101010","000000000000001101","000000000000000101","111111111111110101","111111111111100101","111111111111101101","111111111111011111","111111111111111110","111111111111110100","000000000000101000","000000000000011110","000000000000100010","000000000000001001","000000000000010101","000000000000000110","111111111111110001","000000000000010000","000000000000000011","111111111111100001","000000000000001100","000000000000000001","000000000000010110","111111111111110011","000000000000011010","000000000000000010","000000000000010011","111111111111110100","111111111111101011","111111111111100001","111111111111111101","111111111111110011","111111111111110011","111111111111111001","111111111111111010","111111111111111101","111111111111111100","111111111111100101","111111111111101001","111111111111110101","000000000000100101","111111111111101111","000000000000100101","000000000000000011","111111111111111111","111111111111100101","111111111111110001","111111111111110000","000000000000001000","000000000000001010","111111111111110100","111111111111111110","111111111111110101","000000000000010011","000000000000001011","000000000000010011","111111111111111000","111111111111111001","000000000000010101","000000000000000010","000000000000000011","111111111111011111","111111111111011011","000000000000000001","000000000000010000","000000000000010110","111111111110110010","000000000000011000","000000000000110011","000000000000001011","111111111111110101","000000000000001011","000000000000000001","000000000000000110","111111111111101110","000000000000000100","000000000000001100","111111111111110100","000000000000000010","111111111111100101","000000000000000011","000000000000001100","000000000000010010","000000000000000111","000000000000000010","000000000000001100","000000000000011111","111111111111101011","111111111111100110","111111111111011101","111111111111111011","000000000000010010","000000000000000100","000000000000001000","000000000000010100","000000000000011101","111111111111100101","000000000000000101","111111111110111101","000000000000001110","111111111111110001","000000000000001000","000000000000000110","111111111111110100","000000000000001000","111111111111111100","000000000000000100","000000000000001100","000000000000010010","000000000000000110","111111111111101110","000000000000011011","111111111111101001","000000000000000001","111111111111111110","000000000000001000","000000000000000100","111111111111111110","111111111111111000","000000000000001000","000000000000001011","000000000000010010","000000000000000111","000000000000001000","111111111111101101","000000000000001111","000000000000001001","000000000000001100"),
("000000000000001111","000000000000100010","000000000000001100","111111111111101000","111111111111001010","000000000000001100","111111111111100101","111111111111111001","000000000000000010","000000000000001010","000000000000100000","000000000000010110","000000000000100110","111111111111111110","000000000000010011","111111111111110001","111111111111101110","000000000000001010","000000000000000001","111111111111110011","000000000000001100","000000000000000011","111111111111110100","000000000000010011","000000000000001101","000000000000001001","000000000000100000","111111111111011010","111111111111011100","111111111111101101","000000000000011001","000000000000010001","111111111111110001","000000000000101010","000000000000001110","111111111111111100","000000000000000010","111111111111110011","111111111111111010","111111111111111001","000000000000100010","000000000000010101","000000000000010000","000000000000010001","000000000000011100","111111111111010010","111111111111101110","111111111111110100","000000000000000100","111111111111101001","111111111111101000","000000000000001000","111111111111110010","000000000000010110","111111111111110101","111111111111111000","000000000000000011","111111111111111110","000000000000000110","111111111111110101","000000000000001111","111111111110101010","111111111111011111","111111111111101010","000000000000001011","000000000000100000","111111111111010100","111111111111110010","000000000000111101","000000000000100100","000000000000001101","000000000000000000","111111111111110100","111111111111101101","000000000000000110","111111111111100001","000000000000000000","111111111111110000","111111111111111011","111111111111100110","111111111111110001","111111111111111101","000000000000001010","000000000000010000","111111111111101101","000000000000010000","000000000000011001","111111111111100100","111111111111111010","111111111111100000","000000000000000010","111111111111111000","111111111111110001","111111111111110011","111111111111110000","000000000000001011","111111111111101011","111111111111111111","111111111111110011","000000000000001100","000000000000001011","000000000000001010","000000000000000000","111111111111101111","000000000000100000","111111111111101001","000000000000000100","111111111111101111","000000000000010010","000000000000010000","111111111111110110","000000000000010111","000000000000001110","111111111111110011","000000000000001111","111111111111110101","111111111111111101","000000000000100000","000000000000001111","111111111111101111","000000000000011010","000000000000100110","111111111111111001","000000000000010111","111111111111100110","000000000000001101","000000000000011011","000000000000000100"),
("000000000000001001","000000000000010110","000000000000000011","111111111111110010","111111111110110010","000000000000001011","111111111111100100","111111111111101110","111111111111111001","111111111111111101","000000000000101010","000000000000000011","000000000000010010","000000000000000000","111111111111110111","000000000000001001","111111111111110000","111111111111101010","000000000000010000","000000000000000010","000000000000110010","000000000000000011","111111111111110010","000000000000110010","000000000000001000","000000000000000100","000000000000000100","111111111111100101","111111111111110000","111111111111110011","111111111111111101","000000000000010100","000000000000001011","000000000000001111","000000000000000100","111111111111101100","000000000000001110","000000000000000000","000000000000001110","000000000000100001","000000000000101100","111111111111110011","000000000000011000","000000000000000101","111111111111111110","111111111111011101","111111111111101101","111111111111110110","000000000000010101","111111111111010010","000000000000000100","000000000000001101","111111111111100110","000000000000011001","000000000000001100","111111111111111100","000000000000001100","000000000000000000","000000000000010000","000000000000001011","000000000000100011","111111111110110100","111111111111010111","111111111111101101","111111111111101100","000000000000001100","111111111111111000","111111111111110011","000000000000111101","000000000000011100","111111111111110010","000000000000000000","111111111111111101","000000000000000110","000000000000010100","000000000000000110","111111111111111011","111111111111101101","000000000000000110","111111111111111100","111111111111111010","111111111111110010","000000000000000000","111111111111011000","000000000000000100","111111111111111100","000000000000000000","000000000000000100","000000000000001101","111111111111101100","000000000000000100","111111111111110101","111111111111100101","111111111111110001","111111111111110100","000000000000001011","111111111111101111","000000000000001011","111111111111111110","111111111111111110","111111111111111011","111111111111011110","000000000000001111","111111111111110000","000000000000100010","111111111111101010","111111111111110001","000000000000000111","000000000000001110","000000000000000011","000000000000010010","000000000000001010","000000000000010100","111111111111110001","000000000000001111","111111111111101110","000000000000000010","000000000000001101","000000000000010001","000000000000010001","000000000000010111","000000000000011101","111111111111111000","000000000000010100","000000000000000000","000000000000000000","000000000000001001","000000000000000000"),
("000000000000010000","111111111111111101","000000000000000111","111111111111110010","111111111111000111","000000000000000000","000000000000000000","000000000000011001","000000000000010010","000000000000101101","000000000000110011","000000000000001001","000000000000011001","000000000000000101","111111111111100011","000000000000000010","111111111111011011","000000000000001001","000000000000010111","000000000000001010","000000000001000100","111111111111110111","111111111111111101","000000000000101110","000000000000000000","000000000000000011","111111111111010010","111111111111110110","111111111111101111","111111111111110110","111111111111110111","111111111111111101","111111111111101011","000000000000011111","000000000000000000","111111111111111000","000000000000010110","000000000000100000","111111111111110111","000000000000001011","000000000000011110","111111111111110110","000000000000000110","111111111111111110","000000000000010111","000000000000010110","111111111111110100","111111111111001110","000000000000010100","111111111111100100","000000000000001101","111111111111110110","111111111111100100","000000000000100100","000000000000011110","000000000000001111","000000000000011001","000000000000001000","111111111111111101","000000000000001111","000000000000000010","111111111110001110","111111111111010101","111111111111111100","000000000000010001","111111111111110010","000000000000101001","000000000000000011","000000000000011111","000000000000011101","000000000000000110","000000000000001011","000000000000001111","000000000000010010","000000000000001111","111111111111100101","111111111111110111","111111111111011100","000000000000000000","000000000000000111","000000000000100101","000000000000001000","111111111111111111","111111111110100010","111111111111111011","000000000000011001","111111111111010101","111111111111100001","111111111111101010","000000000000100001","000000000000011110","111111111111110001","111111111111001010","000000000000001000","000000000000000111","111111111111110011","000000000000010110","111111111111111101","000000000000001010","000000000000000011","111111111111111110","111111111110111011","111111111111110101","111111111111110100","000000000000101011","000000000000010010","000000000000100000","000000000000010100","000000000000000111","000000000000001000","000000000000011101","111111111111101111","111111111111111110","111111111111110110","000000000000001100","000000000000001011","111111111111111000","000000000000101111","000000000000000000","000000000000011001","000000000000010110","000000000000001101","111111111111111000","000000000000011110","111111111111111110","111111111111110010","000000000000001100","111111111111111000"),
("000000000000001110","111111111111110111","111111111111111111","111111111111111101","000000000000001101","000000000000010001","111111111111111010","000000000000001100","000000000000001001","000000000000101000","000000000000100011","111111111111010110","000000000000011010","000000000000000000","111111111111110100","000000000000001110","111111111111001001","111111111111110010","000000000000000111","000000000000001110","000000000000110011","111111111111111100","111111111111010100","000000000000010011","000000000000010101","000000000000000101","111111111111001010","111111111111111111","111111111111010111","000000000000010000","000000000000000101","000000000000001101","000000000000001000","000000000000000010","000000000000000110","111111111111101011","000000000000000101","000000000000000000","111111111111100000","000000000000010010","000000000000101001","000000000000000000","000000000000101101","000000000000100111","111111111111110101","000000000000011010","000000000000000101","111111111110111001","000000000000001111","000000000000000000","000000000000000011","000000000000001010","111111111111110010","000000000000100011","000000000000000010","000000000000001111","000000000000000100","000000000000101001","000000000000100000","111111111111111001","111111111111111001","111111111110100111","111111111111100001","111111111111111001","000000000000011011","000000000000000111","000000000000100101","000000000000001000","000000000000101101","000000000000010110","000000000000000001","000000000000100001","000000000000010101","000000000000110000","111111111111110101","000000000000000110","000000000000000001","111111111111011001","111111111111111000","111111111111111010","000000000000000101","111111111111111010","111111111111111011","111111111110110101","111111111111101111","000000000000001110","111111111111010000","111111111111101001","000000000000001110","000000000000101011","000000000000100011","111111111111110111","111111111111011101","000000000000101111","111111111111101110","111111111111111010","000000000000001110","111111111111110001","000000000000100110","111111111111110100","111111111111101111","111111111110111111","000000000000000000","000000000000000011","000000000000010011","111111111111111010","000000000000001011","111111111111110101","111111111111110101","111111111111110011","000000000000011111","000000000000001111","111111111111110111","111111111111111010","111111111111101100","111111111111110101","000000000000000100","000000000000100100","111111111111111001","000000000000011111","111111111111111100","111111111111100010","000000000000010000","000000000000001010","111111111111111101","111111111111110100","000000000000001101","111111111111110101"),
("111111111111111010","111111111111011000","000000000000100001","111111111111100100","000000000000111100","000000000000011000","000000000000000010","000000000000001001","000000000000100000","111111111111110111","000000000000011100","111111111111101000","000000000000011101","000000000000101001","111111111111101111","000000000000010001","111111111111011000","000000000000000001","000000000000010111","111111111111111011","000000000001000110","111111111111101010","111111111111001000","000000000000001011","111111111111111111","000000000000001000","111111111111000110","000000000000010001","111111111111110111","000000000000000100","111111111111110000","111111111111100110","111111111111111011","111111111111101101","000000000000011001","000000000000000011","000000000000000101","000000000000001000","000000000000000110","000000000000000101","111111111111111011","111111111111101011","000000000000010010","000000000000100101","111111111111111001","000000000000101011","111111111111110011","111111111111001010","111111111111110011","000000000000010101","000000000000010000","111111111111100111","000000000000010101","000000000000100110","000000000000101001","000000000000000001","111111111111111000","000000000000010100","000000000000001110","111111111111110000","000000000000000000","111111111111100010","111111111111110010","000000000000000000","000000000000011111","111111111111110111","000000000000100111","111111111111101100","000000000000001000","000000000000000010","111111111111111111","000000000000010100","000000000000011110","000000000000110111","111111111111101011","111111111111111001","111111111111110100","000000000000000100","000000000000000000","111111111111110111","111111111111101111","111111111111100100","111111111111011100","111111111111111000","111111111111110010","000000000000010100","111111111111010111","111111111111110100","000000000000010100","000000000000111000","111111111111011101","111111111111111100","111111111111100110","000000000000110111","000000000000011111","111111111111011111","000000000000011001","000000000000010011","000000000000010100","111111111111011000","000000000000001101","111111111111100110","000000000000000100","000000000000001000","000000000000001111","111111111111111000","000000000000100110","111111111111101001","111111111111111100","111111111111101111","000000000000001000","000000000000001000","111111111111101100","111111111111111101","111111111111110011","000000000000000001","111111111111101100","000000000000100000","000000000000011111","000000000000000001","111111111111111101","111111111111101110","111111111111111010","000000000000001000","000000000000001010","111111111111000111","000000000000010011","000000000000010100"),
("000000000000000011","111111111111011110","000000000000100001","000000000000010000","000000000000111101","111111111111101011","111111111111101011","000000000000000000","000000000000000110","111111111111110011","000000000000000110","000000000000001110","111111111111111111","000000000000010111","111111111111100111","000000000000011101","000000000000010100","111111111111111110","000000000000010000","000000000000011001","000000000000100001","111111111111010011","000000000000000011","111111111111100110","000000000000000110","000000000000000111","000000000000000101","000000000000000100","000000000000011111","000000000000001001","111111111111101101","111111111111110000","111111111111111110","111111111111010100","000000000000001001","000000000000010000","000000000000000111","000000000000010011","111111111111110111","000000000000000111","111111111111100111","111111111111001101","000000000000000111","000000000000010101","000000000000000011","000000000000010011","111111111111101011","111111111111110110","000000000000010000","000000000000010010","000000000000010100","111111111111110000","000000000000000000","000000000000000000","000000000000011111","111111111111111101","111111111111101101","000000000000100100","000000000000100010","111111111111111001","000000000000000100","000000000000010101","000000000000100101","111111111111110000","000000000000000101","000000000000010001","000000000000100010","000000000000000000","111111111111111000","000000000000000101","000000000000010100","000000000000000111","000000000001000011","000000000000110110","111111111111011000","111111111111111101","111111111111101111","000000000000001110","111111111111111110","000000000000010001","000000000000000000","111111111111111000","111111111111110011","000000000000100101","000000000000000101","000000000000010011","111111111111101010","000000000000000010","111111111111111111","000000000000000101","111111111111001111","000000000000000110","000000000000001110","000000000000000000","000000000000011100","111111111111011011","000000000000110101","111111111111111100","111111111111011010","111111111110100001","000000000000001011","000000000000001011","000000000000000000","111111111111110110","000000000000000111","000000000000001000","000000000000000111","111111111111101110","000000000000011001","000000000000001111","000000000000011100","000000000000010101","111111111111110100","000000000000010011","111111111111100111","111111111111111010","000000000000000100","000000000000011011","000000000000001100","000000000000001111","111111111111110100","111111111111111001","111111111111111110","000000000000000010","000000000000010111","111111111111011110","000000000000000111","000000000000000110"),
("111111111111110001","111111111111111101","000000000000011001","000000000000000110","000000000000110110","000000000000000001","111111111111110000","000000000000001110","000000000000000101","111111111111111101","111111111111101110","000000000000001000","000000000000001011","000000000000011011","000000000000000000","000000000000001010","000000000000001010","111111111111110100","000000000000001111","000000000000000111","000000000000110001","111111111111101000","000000000000111011","000000000000000011","000000000000001011","000000000000001000","000000000000010100","000000000000001000","000000000000101111","000000000000000000","000000000000001101","000000000000000111","000000000000001110","111111111110111000","000000000000010100","000000000000000101","111111111111111100","000000000000011010","000000000000010100","000000000000001010","111111111111110010","111111111111000001","000000000000100100","000000000000001101","000000000000000001","111111111111100111","000000000000001000","111111111111100101","000000000000001001","000000000000011011","000000000000001101","000000000000001101","000000000000000001","000000000000000011","000000000000011010","000000000000001100","111111111111111100","000000000000001101","000000000000010101","000000000000001101","000000000000100011","000000000000010111","000000000000110100","000000000000001100","111111111111011010","111111111111111111","000000000000010110","111111111111101001","111111111111111101","000000000000011001","000000000000000100","000000000000011000","000000000000110110","000000000000101101","111111111111011011","111111111111111001","111111111111110001","000000000000010110","000000000000001000","000000000000011000","111111111111110001","000000000000000001","000000000000001011","000000000000110100","000000000000001110","111111111111111110","111111111111100111","111111111111111010","111111111111101010","000000000000000100","111111111111010110","000000000000001111","000000000000101101","111111111111101100","000000000000011100","111111111111100000","000000000000100011","111111111111110101","111111111111100101","111111111111011000","111111111111110010","111111111111101110","000000000000001101","111111111111110011","000000000000010111","111111111111110101","000000000000100111","111111111111110100","000000000000011011","000000000000000000","000000000000000110","000000000000000100","111111111111101001","000000000000010100","111111111111110111","111111111111100111","000000000000000011","000000000000001111","000000000000000010","111111111111111111","111111111111111010","000000000000001110","111111111111100000","000000000000010101","111111111111101001","111111111111010101","111111111111110111","000000000000011101"),
("000000000000000001","111111111111110111","000000000000010110","000000000000100001","111111111111111101","000000000000000000","111111111111110010","111111111111110100","000000000000010111","111111111111101111","000000000000000111","000000000000000101","000000000000000111","000000000000001011","000000000000000110","000000000000010111","000000000000101010","000000000000001100","000000000000000110","000000000000011110","000000000000101000","111111111111111011","000000000000110001","111111111111110110","000000000000001101","000000000000001011","000000000000010000","000000000000001100","000000000000110010","000000000000011001","000000000000000001","111111111111101001","000000000000011011","111111111110111000","111111111111101100","000000000000010111","000000000000011011","000000000000000101","000000000000001111","000000000000011110","000000000000000011","111111111111000010","111111111111110100","000000000000001100","000000000000001100","111111111111111011","111111111111111001","111111111111100001","000000000000001010","000000000000011111","111111111111111100","111111111111111001","000000000000011110","111111111111111001","000000000000011101","000000000000001001","111111111111101100","000000000000011001","000000000000001010","111111111111110001","000000000000000010","000000000000000110","000000000000101110","000000000000010011","111111111111101111","111111111111111010","000000000000101000","111111111111110000","000000000000001010","000000000000101101","111111111111110110","111111111111110101","000000000000111010","000000000000011101","111111111111001001","111111111111010001","111111111111110110","000000000000000000","000000000000000111","000000000000000000","000000000000010111","111111111111111001","000000000000001000","000000000000010001","000000000000010001","000000000000000101","111111111111101000","111111111111101011","111111111111011101","111111111111011001","111111111111100101","111111111111101111","000000000000101110","111111111111010011","000000000000101001","111111111111100000","111111111111101010","111111111111111010","111111111111001011","000000000000010001","000000000000001011","111111111111110110","000000000000000011","000000000000000000","000000000000011011","111111111111111011","000000000000011111","000000000000000010","000000000000101101","111111111111101100","000000000000011100","000000000000010001","111111111111111101","000000000000001010","111111111111110100","000000000000010101","111111111111110010","000000000000000010","000000000000001100","000000000000001101","111111111111111010","000000000000010000","111111111111100001","000000000000011011","111111111111110000","111111111111001000","000000000000001101","000000000000000101"),
("111111111111111010","111111111111111010","000000000000001111","000000000000011000","111111111111011010","111111111111110000","000000000000010110","111111111111111011","111111111111111010","000000000000010100","000000000000000001","111111111111110011","000000000000001000","000000000000011001","111111111111110010","000000000000001001","000000000000100001","000000000000001101","000000000000001011","000000000000011101","111111111111111011","000000000000010011","000000000001000010","111111111111110011","000000000000010011","000000000000000001","000000000000010000","000000000000011101","000000000000100000","000000000000010101","000000000000000101","000000000000001001","000000000000001110","111111111110100100","111111111111110110","000000000000010110","000000000000001000","000000000000001000","000000000000010010","000000000000000011","111111111111110001","111111111110111101","111111111111001000","000000000000001100","000000000000000000","111111111111110010","111111111111101110","111111111111110010","000000000000000101","000000000000110010","000000000000000101","000000000000001011","000000000000011000","111111111111111000","111111111111101011","000000000000001011","000000000000000010","000000000000010111","000000000000011001","111111111111111111","000000000000011100","111111111111100111","000000000000101001","000000000000001001","111111111111101011","000000000000000010","000000000000101110","111111111111101110","111111111111110010","000000000000010011","000000000000010111","000000000000001001","000000000000100011","111111111111110011","111111111111100100","111111111111101011","000000000000000000","000000000000011011","111111111111110100","000000000000000101","000000000000000111","111111111111110110","111111111111111001","111111111111111110","111111111111111000","111111111111101000","111111111111010101","111111111111111101","111111111111011110","111111111111011001","111111111111100011","111111111111110000","000000000000110001","111111111111110010","000000000000010110","111111111111100111","111111111111010111","111111111111110100","111111111111011111","000000000000111111","111111111111111110","111111111111101101","000000000000010100","111111111111111111","000000000000010100","000000000000001000","000000000000010111","000000000000001101","000000000000001001","000000000000000010","000000000000011111","000000000000000101","111111111111110100","000000000000000001","000000000000001001","000000000000001110","111111111111111101","000000000000010011","111111111111111010","111111111111101111","000000000000000010","111111111111110011","111111111111100111","000000000000000010","111111111111101101","111111111111010100","000000000000001111","000000000000000101"),
("111111111111111100","000000000000010101","000000000000010111","111111111111111101","111111111111011111","111111111111110111","000000000000011011","111111111111110000","111111111111110110","000000000000000011","111111111111110111","111111111111110001","111111111111110011","111111111111111101","000000000000001010","111111111111111001","000000000000001111","000000000000010100","000000000000011010","000000000000010011","000000000000000000","000000000000101100","000000000000010011","000000000000010100","000000000000000000","000000000000000100","000000000000100011","000000000000010001","111111111111111101","000000000000000010","111111111111100110","000000000000000100","000000000000010010","111111111110101010","111111111111101111","000000000000010110","000000000000001100","111111111111110110","000000000000010011","000000000000010110","111111111111110101","111111111111001001","111111111110110000","111111111111010110","111111111111110100","111111111111011001","111111111111101101","111111111111101101","000000000000001000","000000000000101010","000000000000010111","000000000000000011","000000000000010101","111111111111001110","000000000000001101","000000000000000101","111111111111011111","000000000000100110","000000000000100011","111111111111110001","111111111111111111","111111111111101000","000000000000001001","111111111111111110","111111111111001000","000000000000010001","000000000000011100","111111111111101001","111111111111111111","000000000000101111","000000000000001000","000000000000011000","000000000000101010","111111111111010001","111111111111100111","111111111111111111","111111111111111001","111111111111111100","000000000000011010","000000000000011110","000000000000001100","000000000000000011","000000000000000111","111111111111110111","000000000000000011","111111111111110000","111111111111011100","111111111111101100","111111111111011110","111111111110111101","000000000000001101","000000000000000001","000000000000100010","000000000000000110","111111111111101011","000000000000000010","111111111110101111","000000000000000011","111111111111110011","000000000001000110","111111111111111111","111111111111101000","000000000000100000","000000000000010010","000000000000010011","000000000000000100","000000000000011001","000000000000011110","111111111111111111","111111111111110100","000000000000011100","111111111111110000","111111111111110001","000000000000000010","000000000000001110","000000000000110001","000000000000001000","000000000000010100","111111111111111100","111111111111101010","111111111111101010","000000000000000100","111111111111010110","000000000000000011","000000000000000111","111111111111100101","000000000000011000","000000000000000110"),
("000000000000101100","111111111111110000","000000000000011101","000000000000001011","111111111111000111","111111111111111111","111111111111111110","111111111111110110","000000000000001000","000000000000001101","000000000000001000","111111111111110100","111111111111101001","111111111111101101","000000000000000000","111111111111101000","000000000000000001","000000000000000101","000000000000000111","000000000000000110","000000000000000101","000000000000100000","000000000000010101","000000000000000111","111111111111100011","000000000000000011","000000000000010111","111111111111110011","111111111111001011","000000000000001001","000000000000000101","000000000000000011","000000000000000001","111111111111001110","000000000000010001","000000000000000000","111111111111111100","111111111111111101","000000000000100110","000000000000011100","111111111111101111","111111111111100010","111111111111000101","111111111111010010","000000000000001001","111111111111100011","111111111111101110","000000000000001011","000000000000100001","000000000000011010","000000000000010100","000000000000000000","000000000000010010","111111111111100100","111111111111100010","000000000000001110","111111111111111110","000000000000000011","000000000000010111","111111111111101010","000000000000011010","111111111111111011","111111111111110011","000000000000001101","111111111111011001","000000000000001001","000000000000010011","111111111111111011","111111111111001011","000000000000100101","000000000000001000","000000000000000101","000000000000101011","111111111110110010","111111111111100000","111111111111111010","111111111111111011","111111111111101110","000000000000000110","000000000000100111","000000000000010001","111111111111111110","111111111111111100","111111111111111001","000000000000001100","111111111111101001","111111111111111011","111111111111110010","111111111111100111","111111111110111001","000000000000010001","000000000000000100","000000000000100001","111111111111111100","111111111111100110","111111111111101010","111111111111000011","111111111111101111","111111111111101011","000000000001010101","000000000000001010","111111111111110011","000000000000000010","111111111111110110","000000000000011100","000000000000010011","000000000000001001","000000000000101000","000000000000000111","111111111111011110","000000000000001101","000000000000000101","000000000000010011","000000000000000011","000000000000101100","000000000000100001","111111111111111001","111111111111111111","000000000000000000","000000000000000101","111111111111101111","111111111111111001","111111111111111000","000000000000001101","000000000000000000","111111111111100001","000000000000000010","000000000000000100"),
("000000000000001011","111111111111110100","000000000000011101","000000000000010100","111111111111010101","111111111111100100","111111111111111110","000000000000000001","111111111111101000","000000000000010100","000000000000000000","111111111111011110","000000000000000110","000000000000001100","111111111111110101","000000000000000000","111111111111011001","000000000000001111","000000000000100101","000000000000010010","000000000000010100","000000000000011111","000000000000000111","111111111111110011","111111111111111000","111111111111110101","000000000000001100","111111111111110101","111111111111010100","000000000000100100","000000000000000000","111111111111111110","000000000000000010","111111111111100001","000000000000001110","111111111111110011","000000000000000010","111111111111111001","000000000000101111","000000000000011000","000000000000000110","111111111111011000","111111111111010001","111111111111011101","000000000000011010","111111111111010011","111111111111110100","111111111111100110","000000000000011110","111111111111111101","000000000000011100","000000000000001110","000000000000010011","111111111111101011","111111111111111110","000000000000010101","111111111111111010","000000000000010010","000000000000010001","111111111111111010","000000000000011111","111111111111111101","111111111111110000","000000000000000010","000000000000000010","111111111111101110","000000000000000001","111111111111100000","111111111111111000","000000000000000001","000000000000010111","000000000000111100","000000000000101101","111111111110101001","111111111111111001","000000000000000001","000000000000000010","000000000000001011","000000000000000111","000000000000100100","111111111111110001","111111111111111111","111111111111101111","000000000000001100","000000000000000100","111111111111011001","000000000000000001","111111111111111000","111111111111101110","111111111111000011","111111111111111101","111111111111110111","000000000000001000","111111111111101001","111111111111101111","111111111111110111","111111111111010001","111111111111111011","000000000000010001","000000000000110011","111111111111100001","111111111111110010","000000000000001110","111111111111110100","000000000000011100","000000000000011111","111111111111111010","000000000000000001","000000000000010010","111111111111011101","000000000000000000","111111111111111000","111111111111110001","000000000000011001","000000000000111100","000000000000000110","000000000000000000","000000000000010110","000000000000001011","000000000000010011","111111111111111010","000000000000000111","111111111111111010","111111111111110101","111111111111111100","111111111111000001","000000000000011100","111111111111110100"),
("000000000000000001","111111111111110100","000000000000001100","000000000000001011","111111111111011101","111111111111110101","000000000000000000","111111111111110001","000000000000000111","000000000000010101","000000000000011011","111111111111101000","111111111111110111","111111111111011100","111111111111101010","000000000000011100","111111111111011111","000000000000101010","000000000000001010","111111111111111101","000000000000001011","000000000000110011","111111111111110010","000000000000011011","111111111111110111","000000000000000001","000000000000100110","111111111111100011","111111111111000111","000000000000010111","111111111111111110","111111111111101111","000000000000011011","111111111111110100","111111111111111101","111111111111100110","111111111111110101","111111111111101011","000000000000001000","000000000000000110","000000000000000011","111111111111010000","111111111111101000","111111111111011111","000000000000011001","111111111111100001","111111111111110110","111111111111010000","000000000000011000","000000000000001010","000000000000010001","000000000000011101","000000000000001110","111111111111001011","000000000000000011","000000000000100001","111111111111110111","000000000000010001","111111111111111111","111111111111110010","000000000000000101","111111111111111010","111111111111101101","111111111111111011","111111111111110101","111111111111110111","000000000000010111","111111111111111011","111111111111111010","000000000000001100","000000000000000000","000000000000010101","000000000000100101","111111111110011111","111111111111010011","111111111111101001","111111111111110010","000000000000001100","111111111111111001","000000000000011010","111111111111101110","000000000000001111","111111111111111101","111111111111110110","000000000000010011","111111111111111000","000000000000000100","111111111111011011","111111111111101101","111111111111100110","000000000000000001","111111111111111000","000000000000001100","000000000000010000","111111111111100001","111111111111011000","111111111111011111","000000000000000001","111111111111111000","000000000000000100","111111111111100110","111111111111111110","000000000000001011","000000000000010001","000000000000100000","000000000000001111","111111111111110011","000000000000000101","111111111111110111","111111111111101100","000000000000001101","111111111111110110","000000000000001101","000000000000001100","000000000001000001","000000000000000001","111111111111110010","000000000000001110","000000000000011101","000000000000001000","111111111111110101","111111111111110101","111111111111100011","000000000000001010","111111111111110100","111111111110111111","000000000000001110","111111111111110011"),
("000000000000110001","000000000000010000","000000000000011001","111111111111010010","111111111110110011","111111111111101101","111111111111110111","111111111111101010","111111111111101101","000000000000001000","111111111111101110","000000000000001110","111111111111111101","111111111111110010","111111111111101000","000000000000000110","111111111111011101","000000000000001000","111111111111111010","111111111111110000","000000000000110001","000000000000101001","000000000000000100","000000000000010100","000000000000010101","111111111111110011","000000000000011011","111111111111010101","111111111111010110","000000000000011001","000000000000010011","111111111111100000","000000000000000110","111111111111101000","000000000000110001","111111111111101000","000000000000101001","111111111111111010","000000000000110010","000000000000011000","000000000000101011","000000000000000010","111111111111110100","111111111111001101","000000000000010111","111111111111110110","111111111111101110","111111111111101011","000000000000011011","111111111111000011","000000000000010101","000000000000110000","000000000000111001","111111111111100000","111111111111111100","000000000000000001","000000000000011010","111111111111110100","000000000000000101","111111111111111111","000000000000010001","111111111111011101","111111111110110111","111111111111100001","111111111111110110","000000000000110111","000000000000011010","000000000000001000","111111111111100110","000000000000110100","111111111111111101","000000000000000000","000000000000001100","111111111111010011","111111111110111011","111111111111111110","000000000000011001","111111111111010111","000000000000000001","111111111111111111","000000000000010000","000000000000000100","111111111111100001","111111111111010100","000000000000100010","111111111111101010","000000000000001000","111111111111100001","000000000000000000","111111111111101100","000000000000011101","000000000000000111","000000000000110111","111111111111101100","111111111111111001","111111111111011100","111111111111110000","111111111111111101","000000000000001111","111111111111110110","000000000000000111","000000000000000111","111111111111101110","000000000000001000","000000000000110011","111111111111111010","000000000000000111","000000000000001010","111111111111110011","000000000000010101","000000000000010111","111111111111111100","000000000000010100","000000000000000000","000000000000001101","111111111111101110","111111111111100011","000000000000010010","000000000000101010","111111111111110010","111111111111111100","000000000000110100","111111111111110010","000000000000001111","111111111111100110","111111111111111110","000000000000000010","111111111111111101"),
("000000000000001100","000000000000001011","000000000000100010","000000000000001011","111111111111011110","111111111111101010","000000000000000101","000000000000001110","000000000000001110","000000000000001001","111111111111110010","000000000000010110","111111111111110110","111111111111000110","111111111111100100","000000000000001010","111111111111100001","000000000000111010","000000000000100100","111111111111111111","000000000000001101","111111111111110100","111111111111010000","000000000000001010","000000000000011100","000000000000000011","000000000000101011","111111111111011101","111111111111101100","000000000000101110","000000000000100110","111111111111010100","111111111111110110","111111111111110110","000000000000100101","111111111111111110","000000000000000000","000000000000010011","000000000000100101","000000000000010110","000000000000010101","000000000000100000","000000000000001000","111111111111101110","000000000000101101","111111111111110000","111111111111111001","000000000000011100","000000000000110100","111111111111010001","000000000000001101","000000000000100010","000000000000001101","111111111111101100","111111111111111101","000000000000000011","000000000000110111","111111111111101111","111111111111101100","000000000000001001","000000000000100001","111111111111111111","111111111111101111","111111111111101111","111111111111010101","000000000000111000","000000000000010100","000000000000000101","111111111111110101","000000000000010110","000000000000000000","000000000000000100","000000000000001101","111111111111100001","111111111111100101","000000000000001110","000000000000011010","111111111111100001","111111111111101000","000000000000001110","000000000000000110","000000000000011010","111111111111001011","111111111111100101","000000000000101000","111111111110111101","111111111111111000","000000000000000010","000000000000001100","111111111111100101","000000000000010110","000000000000001110","000000000000001110","111111111111010101","111111111111100011","111111111111111111","000000000000000010","111111111111111000","000000000000100101","111111111111111001","000000000000001101","111111111111111100","111111111111011001","000000000000101100","000000000000111100","000000000000001111","111111111111111100","000000000000000001","111111111111100000","111111111111101001","000000000000001000","111111111111110010","000000000000101101","000000000000001011","000000000000110011","111111111110111001","111111111111011100","000000000000001100","000000000000011011","000000000000000000","111111111111101100","111111111111111111","111111111111110011","111111111111110110","111111111111011001","111111111111101000","000000000000100001","000000000000011010"),
("111111111111111010","111111111111001111","111111111111101001","000000000000001110","111111111111001010","111111111111111111","111111111111110010","111111111111111101","000000000000010001","111111111111001000","111111111111111010","000000000000001101","000000000000100001","111111111111100100","000000000000000001","111111111111011101","111111111111011001","000000000000110000","000000000000101000","111111111111101001","000000000000011100","111111111111010101","111111111111010001","111111111111101111","000000000000010111","111111111111111110","000000000000100100","111111111111011111","111111111111110111","111111111111110100","000000000000011011","111111111111100101","111111111111110101","111111111111101100","000000000000111000","111111111111111110","111111111111110000","000000000000100001","000000000000011111","000000000000001000","000000000000011110","000000000000110100","000000000000000110","111111111111011011","000000000000101011","111111111111110000","000000000000001000","111111111111110001","000000000000111101","111111111111111111","111111111111100111","000000000000001000","000000000000000110","000000000000001001","111111111111011111","000000000000011100","000000000000000110","111111111111101101","111111111111101001","111111111111110010","000000000000001111","000000000000010001","111111111111100000","111111111111101111","111111111111100110","000000000000000011","111111111111110111","111111111111111011","000000000000011010","000000000000001101","111111111111110101","000000000000011011","000000000000000100","111111111111101100","111111111111111111","000000000000000100","000000000000010101","111111111111100011","111111111111110111","000000000000010010","111111111111101111","000000000000010011","111111111111101010","000000000000000000","000000000000001111","111111111111011001","000000000000011001","000000000000000100","111111111111100101","111111111111110010","111111111111101110","111111111111111000","000000000000010001","111111111111011000","000000000000010111","111111111111101110","111111111111101110","111111111111111111","000000000000000000","000000000000001000","000000000000000001","000000000000001010","111111111111010001","111111111111111000","000000000000011111","111111111111111100","111111111111111010","000000000000010100","111111111111111100","111111111111101000","000000000000000111","111111111111101110","000000000000000010","000000000000011110","000000000000100001","111111111111011111","111111111111111110","111111111111100101","111111111111111101","111111111111100101","000000000000000100","000000000000000111","111111111111111100","111111111111001000","111111111111111100","111111111111111000","000000000000100000","000000000000001111"),
("111111111111011101","111111111111101001","000000000000011100","111111111111101001","000000000000000101","111111111111101000","000000000000000010","111111111111111111","111111111111110101","111111111111110110","111111111111101011","111111111111111100","000000000000001000","000000000000100000","000000000000001100","000000000000011111","111111111111010001","111111111111101100","000000000000101001","111111111111111001","000000000000101100","111111111111101101","111111111111111111","111111111111111011","000000000000010100","111111111111100011","111111111111101000","000000000000000001","000000000000000010","000000000000000000","111111111111100100","000000000000001011","111111111111101000","000000000000000011","000000000000001011","111111111111101011","000000000000001010","111111111111110101","111111111111101010","000000000000000100","000000000000011110","000000000000100101","000000000000101001","000000000000000000","111111111111111100","111111111111110100","111111111111111101","111111111111011101","000000000000101010","111111111111111000","111111111111110101","111111111111110001","000000000000100011","000000000000001111","000000000000010001","000000000000001100","111111111111100111","111111111111111010","000000000000101010","111111111111111101","111111111111110100","000000000000001011","000000000000000101","111111111111100001","000000000000001010","000000000000100001","000000000000000000","111111111111101110","000000000000110011","000000000000000001","111111111111111001","000000000000001111","000000000000001111","111111111111101100","111111111111110000","111111111111110100","111111111111100010","111111111111100011","000000000000011111","111111111111111100","111111111111011011","111111111111101010","000000000000000011","000000000000010001","111111111111011001","000000000000100101","000000000000001111","000000000000000000","111111111111010010","111111111111101100","111111111111110101","111111111111111011","000000000000001001","111111111111101101","000000000000010000","111111111111110101","111111111111111000","111111111111110110","000000000000001100","000000000000110101","111111111111100101","111111111111100011","000000000000000000","111111111111110011","111111111111100101","111111111111101000","111111111111111000","000000000000010000","000000000000000000","111111111111110101","111111111111111101","111111111111111001","111111111111100001","111111111111110010","000000000000000110","111111111111110111","111111111111100011","000000000000010001","111111111111100001","000000000000001001","000000000000010000","111111111111010110","000000000000001001","111111111111010110","000000000000011101","111111111111100010","000000000000010110","000000000000100100"),
("000000000000000101","111111111111110011","000000000000010011","111111111111101100","000000000000000100","111111111111101100","000000000000001001","000000000000000101","000000000000010110","000000000000010100","000000000000000011","000000000000000011","000000000000010101","000000000000010010","000000000000000100","111111111111111010","000000000000000000","111111111111111100","000000000000010110","000000000000011110","000000000000011110","111111111111110000","111111111111110100","111111111111111111","000000000000001100","111111111111110101","111111111111110000","111111111111110111","000000000000000000","000000000000000010","000000000000001000","111111111111111010","111111111111110110","111111111111110000","111111111111111000","111111111111101100","000000000000011110","111111111111110101","111111111111110010","000000000000001000","000000000000000100","000000000000001000","000000000000010110","111111111111111000","111111111111110110","000000000000011000","111111111111111111","000000000000010000","000000000000001001","000000000000000111","111111111111101101","111111111111101110","000000000000010011","000000000000000011","000000000000011101","000000000000001000","000000000000000010","000000000000011011","000000000000010110","111111111111101111","000000000000001111","111111111111111010","000000000000001001","111111111111101010","000000000000000110","000000000000001111","000000000000001000","111111111111111011","111111111111111001","111111111111110111","111111111111111111","111111111111111101","000000000000001000","000000000000010010","000000000000000001","111111111111111100","000000000000000000","000000000000001001","000000000000001111","000000000000001111","111111111111101101","111111111111111110","111111111111101100","111111111111110000","111111111111111010","000000000000011101","000000000000010100","000000000000001011","000000000000000110","111111111111110110","000000000000011000","000000000000000110","000000000000100011","111111111111111100","000000000000011110","111111111111111000","111111111111111100","111111111111111110","111111111111111101","000000000000000100","111111111111101011","000000000000001011","111111111111110011","111111111111110111","111111111111111110","111111111111101110","000000000000001100","000000000000000100","111111111111101101","000000000000010100","000000000000010011","000000000000000000","111111111111110110","000000000000000001","000000000000010110","000000000000001011","111111111111101110","111111111111111100","111111111111101110","000000000000010101","000000000000001010","000000000000000101","000000000000011010","000000000000011001","000000000000001000","000000000000001000","111111111111111111","111111111111111001"),
("000000000000010110","000000000000000111","000000000000000011","111111111111101110","000000000000011101","000000000000000110","111111111111100011","111111111111011100","111111111111111101","111111111111111010","000000000000000101","111111111111110100","111111111111111001","000000000000001010","000000000000001111","111111111111110001","111111111111110101","000000000000000010","111111111111111001","111111111111111011","000000000000011100","000000000000010100","000000000000011001","111111111111110010","000000000000000011","000000000000001010","000000000000000011","111111111111111110","111111111111110101","000000000000001001","111111111111111001","000000000000011101","000000000000000000","000000000000000010","000000000000000011","111111111111100100","111111111111110111","000000000000001101","000000000000001100","111111111111111111","000000000000000111","000000000000001001","111111111111110111","000000000000001100","111111111111101011","000000000000001000","000000000000001111","111111111111110101","111111111111111000","111111111111110111","000000000000001000","000000000000001101","111111111111110101","000000000000001011","111111111111111000","111111111111110100","000000000000000011","000000000000010111","000000000000001100","111111111111110111","111111111111111010","111111111111111111","000000000000000111","111111111111111001","111111111111111111","000000000000010101","111111111111110111","111111111111101011","111111111111111111","000000000000001000","111111111111100101","000000000000010111","111111111111110111","000000000000000000","111111111111110111","111111111111101100","111111111111110101","111111111111101100","000000000000001001","000000000000001010","111111111111111101","111111111111101101","111111111111111111","000000000000010000","111111111111111111","000000000000000000","000000000000010111","000000000000000101","111111111111100111","111111111111111001","111111111111111011","111111111111110111","000000000000000111","000000000000001100","111111111111111101","111111111111110001","000000000000001000","111111111111110110","000000000000001110","000000000000001010","111111111111111100","111111111111101000","111111111111110010","111111111111111111","111111111111111100","111111111111101011","111111111111101101","000000000000001111","111111111111110011","111111111111111101","111111111111111000","000000000000001010","000000000000000110","000000000000010111","111111111111101110","111111111111110011","111111111111110100","000000000000011001","000000000000000011","000000000000010011","000000000000000101","111111111111111000","000000000000000101","000000000000000100","000000000000011000","111111111111111111","000000000000001101","111111111111110100"),
("111111111111100100","000000000000000000","000000000000010100","111111111111100000","000000000000001000","111111111111100000","111111111111110101","111111111111010010","111111111111110101","000000000000100011","111111111111110010","000000000000001011","000000000000010111","000000000000010111","111111111111111010","111111111111111010","000000000000001011","111111111111111111","000000000000010100","000000000000001101","111111111111110011","000000000000001011","000000000000100111","111111111111110010","111111111111110111","111111111111110001","111111111111111011","111111111111101010","000000000000000100","000000000000010100","111111111111011111","111111111111101110","111111111111111001","111111111111100100","111111111111111001","000000000000000111","000000000000000111","000000000000001001","111111111111110001","000000000000001101","000000000000001101","111111111111111010","000000000000001001","111111111111111110","111111111111100111","111111111111111101","000000000000010101","111111111111111111","000000000000000101","000000000000000000","000000000000000101","000000000000000100","000000000000000100","111111111111100010","000000000000000111","111111111111111000","111111111111101101","000000000000011011","000000000000000111","000000000000000001","000000000000010100","000000000000000111","111111111111100000","000000000000001100","111111111111101111","000000000000100101","000000000000010111","111111111111111100","000000000000010001","000000000000001011","111111111111101110","000000000000010001","111111111111100001","000000000000010010","111111111111010100","111111111111101001","000000000000000000","111111111111100100","111111111111111010","000000000000011011","111111111111111100","111111111111011010","111111111111100101","000000000000011000","111111111111101010","000000000000010110","000000000000011010","000000000000001000","111111111111101010","000000000000010011","111111111111110110","111111111111110101","111111111111101110","000000000000000011","000000000000000000","111111111111100000","111111111111111001","111111111111111010","111111111111110101","111111111111110110","111111111111111011","111111111111101001","111111111111110101","000000000000011001","000000000000000000","111111111111111111","000000000000000011","000000000000011100","111111111111110111","000000000000100010","000000000000000100","111111111111110011","111111111111111110","000000000000001101","000000000000001111","111111111111101100","111111111111101000","000000000000011111","111111111111100010","111111111111101101","000000000000010110","000000000000010000","000000000000001110","111111111111110101","000000000000100001","111111111111101000","000000000000001001","111111111111111111"),
("111111111111011010","000000000000001001","000000000000001010","000000000000000111","111111111111110100","111111111111101111","000000000000000000","111111111111101000","000000000000001010","000000000000010001","000000000000000111","111111111111111101","111111111111111110","000000000000001101","000000000000000000","000000000000001111","000000000000001011","000000000000000000","000000000000001010","000000000000000110","111111111111111010","000000000000001101","000000000000000100","000000000000000010","111111111111101010","111111111111110000","111111111111111111","000000000000000010","000000000000100011","111111111111110110","111111111111100111","000000000000000110","000000000000010101","111111111111110000","111111111111110010","111111111111111101","111111111111110001","000000000000011101","111111111111110100","111111111111111100","111111111111110000","111111111111100010","000000000000011001","000000000000000100","111111111111110111","000000000000001101","000000000000011001","111111111111000100","000000000000010001","000000000000010111","000000000000001101","000000000000010001","000000000000010000","000000000000010001","000000000000101010","000000000000000111","111111111111111011","000000000000000111","111111111111111111","000000000000000110","000000000000000110","111111111111100011","111111111111100110","111111111111110111","111111111111111111","111111111111011111","111111111111101110","000000000000001100","000000000000001010","111111111111101101","000000000000001111","000000000000100101","000000000000000000","000000000000101000","000000000000001000","111111111111110100","111111111111110101","000000000000011011","111111111111111110","000000000000011011","111111111111010111","000000000000000101","000000000000000100","000000000000010011","000000000000001010","000000000000000011","111111111111110011","000000000000000101","000000000000000110","000000000000001001","111111111111100111","111111111111010000","111111111111111001","000000000000001001","111111111111110011","111111111111101000","111111111111111011","111111111111111010","000000000000000111","000000000000000100","000000000000000010","111111111111010110","111111111111101011","111111111111110001","111111111111110100","000000000000010010","000000000000000001","111111111111111110","111111111111111111","111111111111011110","111111111111110010","000000000000010101","111111111111110111","000000000000011001","000000000000101000","000000000000001111","000000000000010010","000000000000001000","111111111111100001","000000000000010111","000000000000000101","111111111111100001","000000000000010010","000000000000001110","111111111111100110","111111111111010011","000000000000000010","000000000000000100"),
("111111111111101011","111111111111110111","000000000000010000","111111111111101101","111111111111110101","111111111111110001","111111111111101100","000000000000010110","000000000000000000","111111111111110010","000000000000001010","000000000000100011","111111111111101100","111111111111110001","000000000000001000","111111111111111010","111111111111010111","000000000000011101","000000000000001010","111111111111100001","111111111111111100","000000000000101100","111111111111100101","000000000000000100","000000000000001011","111111111111111110","000000000000011001","111111111111101101","000000000000011000","111111111111111001","111111111111100111","000000000000000010","111111111111100110","111111111111101101","111111111111110100","000000000000001001","000000000000000010","000000000000100011","000000000000000011","000000000000001011","000000000000100111","000000000000000000","000000000000100101","000000000000001101","111111111111110011","111111111111110111","000000000000010110","111111111111011111","000000000000010100","000000000000001100","000000000000000000","111111111111110110","000000000000000011","000000000000011111","111111111111111000","111111111111111011","111111111111101001","000000000000000101","111111111111111100","111111111111111110","000000000000001001","111111111111100001","111111111111100100","000000000000000000","111111111111111101","000000000000000101","111111111111111000","111111111111111011","000000000000001101","000000000000000001","111111111111110111","000000000000001111","000000000000000011","000000000000010100","000000000000000001","111111111111110000","111111111111101111","111111111111101010","111111111111110111","111111111111011010","000000000000000101","000000000000000101","111111111111100100","111111111111111010","111111111111111010","111111111111111110","000000000000000000","000000000000001000","111111111111001111","000000000000001100","111111111111110011","111111111111100010","000000000000100111","111111111111101101","111111111111110100","111111111111110000","111111111111010011","000000000000000000","111111111111101101","000000000000001000","111111111111110000","111111111111110100","111111111111110100","000000000000001011","000000000000010011","111111111111110010","000000000000001001","111111111111111111","000000000000000000","000000000000000011","000000000000001001","111111111111111000","000000000000010111","000000000000010000","000000000000011001","000000000000001010","111111111111101111","000000000000100000","111111111111101011","111111111111110101","000000000000000000","111111111111110110","111111111111110100","000000000000101100","111111111111100010","111111111111011001","111111111111101100","111111111111101000"),
("111111111111010011","111111111111111001","111111111111111011","111111111111110110","000000000000000101","111111111111111110","000000000000010100","000000000000101000","000000000000011000","111111111111110111","000000000000101100","111111111111111001","000000000000001000","111111111111101000","000000000000000000","000000000000000001","111111111111101111","111111111111111010","111111111111110110","000000000000000110","000000000000000110","000000000000001101","000000000000001101","111111111111110110","111111111111110001","000000000000010101","111111111111110100","000000000000010010","111111111111110110","111111111111100111","000000000000001000","000000000000000110","000000000000100010","111111111111001001","111111111111110110","000000000000001000","000000000000000100","111111111111111010","111111111111111100","111111111111101101","111111111111111100","111111111111100001","000000000000101111","000000000000001010","000000000000001110","111111111111110101","000000000000001101","000000000000000001","111111111111110100","000000000000000101","111111111111110101","000000000000000100","111111111111111010","000000000000101001","000000000000010011","000000000000011000","111111111111100101","000000000000000101","111111111111111001","000000000000000111","111111111111100010","111111111111100100","000000000000000101","111111111111110010","111111111111010100","000000000000100000","111111111111101001","000000000000000000","000000000000011011","111111111111111101","000000000000001000","111111111111110010","000000000000000101","000000000000000110","111111111111110110","000000000000001110","000000000000000010","111111111111100101","000000000000001100","111111111111011111","111111111111100001","000000000000010000","111111111111100111","111111111111010101","000000000000000111","000000000000010100","000000000000001110","111111111111111000","111111111111110100","111111111111101000","111111111111001011","111111111111111101","000000000000000101","111111111111100001","000000000000000011","111111111111111100","111111111111101110","000000000000011000","111111111111011000","000000000000011110","111111111111111011","111111111111101110","111111111111100111","111111111111110100","111111111111100110","000000000000011000","000000000000010101","000000000000010000","111111111111111001","111111111111111000","000000000000000000","000000000000110110","111111111111110110","000000000000001010","000000000000000110","111111111111110010","111111111111110011","000000000000011110","111111111111011001","111111111111111010","000000000000010100","111111111111110010","000000000000000000","000000000000011100","111111111111111001","000000000000000001","000000000000000001","000000000000001010"),
("111111111111010111","000000000000011111","111111111111111101","111111111111101010","111111111111101000","111111111111100001","000000000000100110","000000000000000010","000000000000001001","111111111111101100","000000000000101010","000000000000000110","111111111111111001","111111111111110001","000000000000001110","111111111111101001","111111111111010111","000000000000000001","111111111111110111","000000000000000011","111111111111111110","000000000000010111","111111111111101101","111111111111011011","000000000000000011","111111111111111011","111111111111101110","000000000000001101","111111111111100110","111111111111110000","111111111111110011","111111111111110100","000000000000000000","111111111111100100","111111111111101100","111111111111111111","111111111111111111","000000000000001010","111111111111010110","111111111111110001","000000000000010110","111111111111111000","000000000000100011","000000000000010000","111111111111111010","111111111111101100","111111111111110111","111111111111100111","111111111111110111","000000000000010001","111111111111011011","111111111111110001","000000000000011010","000000000000101001","000000000000010001","000000000000011101","111111111111100101","000000000000011000","000000000000001001","000000000000000000","111111111111111001","111111111111000110","111111111111110010","000000000000001010","111111111110100010","111111111111111111","111111111111011100","111111111111111110","000000000000100011","111111111111111010","000000000000010011","000000000000000101","000000000000000001","000000000000011110","000000000000001011","000000000000010001","111111111111111100","000000000000000010","000000000000001111","111111111111101101","111111111111110100","000000000000001000","111111111111101110","111111111111001101","111111111111110011","111111111111110001","111111111111111001","111111111111101111","000000000000000000","111111111111101110","111111111111011010","000000000000000110","000000000000011000","000000000000001000","000000000000001001","111111111111100100","111111111111001100","000000000000101001","111111111111110001","000000000000000100","000000000000000010","111111111111110010","111111111111010001","111111111111111110","111111111111101111","000000000000010110","000000000000000110","000000000000001100","111111111111111100","111111111111110101","000000000000100011","000000000000010110","111111111111101101","000000000000000110","000000000000101101","111111111111100111","000000000000010011","000000000000100011","111111111111010110","111111111111111110","000000000000010010","111111111111100100","000000000000000101","000000000000110010","111111111111110100","000000000000011001","111111111111111001","111111111111110110"),
("111111111111001011","000000000000011100","111111111111111111","111111111111111000","111111111111110110","111111111111110011","000000000000011110","111111111111011110","000000000000001111","111111111111011101","000000000000111100","000000000000010101","111111111111111110","111111111111101001","000000000000100001","111111111111100100","111111111111011111","111111111111110011","000000000000011000","111111111111010100","000000000000010001","111111111111110111","111111111111101110","111111111111011111","111111111111110001","000000000000000001","000000000000010000","111111111111111100","111111111111111110","111111111111110011","111111111111111100","000000000000010100","111111111111111010","111111111111011010","000000000000001111","111111111111111011","111111111111111101","111111111111111011","000000000000000011","111111111111110010","000000000000001111","111111111111011111","000000000000101101","000000000000001101","000000000000000111","000000000000000100","000000000000100110","111111111111111110","111111111111111010","111111111111111110","111111111111011111","111111111111111100","000000000000001011","000000000000101101","111111111111101110","111111111111111011","000000000000000001","000000000000001100","000000000000100000","000000000000000001","000000000000010010","111111111111000011","111111111111011000","000000000000001110","111111111111100111","000000000000010000","111111111111100011","111111111111111001","000000000000011000","000000000000010111","000000000000000110","000000000000001001","111111111111101000","000000000000010000","000000000000001010","000000000000001110","111111111111111100","000000000000000010","111111111111111100","111111111111011010","000000000000001110","111111111111111011","111111111111101001","111111111111101101","000000000000000010","111111111111111010","000000000000000110","111111111111100011","111111111111111010","111111111111000111","111111111111101010","111111111111111101","000000000000001000","111111111111111100","000000000000010011","111111111111101001","111111111111100000","000000000000010010","000000000000010001","000000000000010000","000000000000001011","000000000000010011","111111111111111110","000000000000000111","111111111111010100","000000000000011001","000000000000000000","000000000000000010","000000000000000001","111111111111110010","000000000000000000","000000000000011100","111111111111111110","000000000000000010","000000000000000100","111111111111100101","111111111111110000","000000000000010000","111111111111100101","111111111111111101","111111111111111000","111111111111100001","111111111111111101","000000000000001100","111111111111110011","000000000000101011","111111111111111011","000000000000001100"),
("111111111111100100","000000000000000110","000000000000010001","111111111111110001","000000000000101000","111111111111111110","000000000000001100","000000000000000100","111111111111100111","111111111111100011","000000000000011001","000000000000010101","000000000000010101","000000000000001100","111111111111111110","000000000000001000","111111111111100100","000000000000000000","000000000000000100","111111111111110110","111111111111110111","000000000000011000","000000000000010001","111111111111000001","111111111111111010","111111111111101110","000000000000010010","111111111111110001","111111111111110000","111111111111100100","000000000000000101","000000000000010000","111111111111110111","000000000000000110","000000000000001101","000000000000001110","000000000000000010","111111111111101110","000000000000001001","111111111111111000","000000000000011000","111111111111111001","000000000000001101","111111111111110010","111111111111111101","111111111111011011","000000000000000000","111111111111111100","000000000000001111","000000000000000100","000000000000000000","111111111111110100","000000000000010000","000000000000101100","000000000000000010","000000000000000000","111111111111110101","000000000000000001","000000000000011000","111111111111110110","111111111111101101","111111111110110111","111111111111010101","111111111111110101","111111111111110100","000000000000001111","111111111111010100","000000000000010011","000000000000100100","111111111111111110","111111111111111001","111111111111111000","111111111111100000","111111111111110111","111111111111111111","000000000000001101","000000000000010011","000000000000000001","000000000000010011","111111111111100101","000000000000000000","000000000000010001","111111111111111101","111111111111111111","111111111111101110","000000000000000000","000000000000001011","111111111111101010","000000000000001000","111111111111001011","111111111111110111","111111111111111110","000000000000100001","111111111111111010","000000000000000101","000000000000000101","111111111111101001","000000000000001001","111111111111110011","000000000000001101","111111111111111101","000000000000110010","111111111111101111","111111111111111000","111111111111011100","111111111111110001","000000000000001100","000000000000000101","000000000000010001","000000000000000111","000000000000000101","000000000000000110","000000000000000000","000000000000000101","000000000000011111","111111111111110100","111111111111101100","000000000000001011","000000000000010000","111111111111111011","000000000000010011","111111111111100101","000000000000000101","000000000000011100","111111111111110011","000000000000011111","000000000000001001","000000000000000110"),
("111111111111111000","000000000000101111","000000000000100001","111111111111110010","000000000000110000","000000000000000010","000000000000000110","111111111111100110","111111111111101111","111111111111111101","000000000000011111","000000000000011000","000000000000001011","111111111111111000","111111111111111010","111111111111101101","111111111111011110","111111111111101001","000000000000000000","111111111111101100","000000000000011101","000000000000001001","000000000000010000","111111111111010010","000000000000010100","111111111111110101","111111111111111110","111111111111100111","111111111111110011","111111111111011111","111111111111110101","000000000000000001","111111111111101101","000000000000000111","000000000000010011","111111111111110111","111111111111111000","111111111111111000","000000000000001001","111111111111111001","000000000000101100","000000000000001100","000000000000011100","000000000000000011","000000000000001110","111111111111001110","111111111111111001","111111111111111111","000000000000010100","000000000000000100","000000000000000001","000000000000000100","000000000000011001","000000000000011111","000000000000000010","111111111111111111","111111111111110100","000000000000000111","111111111111111101","000000000000000100","000000000000000000","111111111110011101","111111111110111010","111111111111110100","111111111111111100","000000000000000011","111111111111001100","000000000000001101","000000000000101101","111111111111111101","111111111111110100","000000000000010001","111111111111100011","000000000000010010","111111111111101111","111111111111110100","000000000000001101","111111111111101011","111111111111111100","111111111111111010","000000000000001010","000000000000000001","111111111111101000","000000000000010010","111111111111110100","000000000000000010","000000000000011000","111111111111110101","111111111111110011","111111111111000011","111111111111111001","000000000000011000","000000000000111001","111111111111100001","000000000000100011","000000000000010111","111111111111011101","000000000000010101","111111111111011001","000000000000011110","111111111111110010","000000000001000000","111111111111111000","000000000000001110","111111111111110111","000000000000000101","111111111111111000","111111111111111100","000000000000000110","000000000000001111","000000000000001011","000000000000010000","111111111111111001","111111111111110110","000000000000001010","000000000000001110","000000000000000011","000000000000001110","000000000000001001","111111111111111100","000000000000010110","000000000000000000","111111111111101010","000000000000010001","111111111111011110","000000000000001001","000000000000000001","000000000000001100"),
("000000000000100011","000000000000101110","000000000000010100","111111111111110110","111111111111111101","111111111111101000","111111111111111100","000000000000000000","111111111111110001","000000000000001010","000000000000111101","000000000000011100","000000000000011000","000000000000010101","111111111111110001","000000000000000111","111111111111001111","111111111111101000","000000000000001011","111111111111101110","000000000000010011","000000000000100010","111111111111101000","000000000000000110","000000000000100011","000000000000000101","000000000000100101","111111111111101100","111111111111111000","111111111111010110","000000000000010011","000000000000001010","111111111111101001","111111111111111101","111111111111111000","000000000000001001","000000000000001100","111111111111100111","111111111111111011","000000000000011010","000000000000011011","111111111111111000","000000000000001010","111111111111110110","111111111111111011","111111111111010110","111111111111111011","000000000000001111","000000000000000111","111111111111111000","111111111111110110","000000000000001011","111111111111111011","000000000000100011","111111111111111000","000000000000010111","000000000000010111","111111111111110010","000000000000010011","000000000000000110","000000000000001000","111111111110001111","111111111110100001","000000000000000000","000000000000011000","000000000000011010","111111111110111010","000000000000000010","000000000000001111","000000000000011011","000000000000000101","111111111111111100","111111111111101011","000000000000000000","000000000000001000","111111111111101000","000000000000010011","111111111111110011","111111111111101110","000000000000000000","000000000000001001","000000000000001000","000000000000000000","111111111111111101","111111111111101111","111111111111111001","000000000000001110","111111111111100101","000000000000001110","111111111111001001","000000000000001110","000000000000011001","000000000000001010","111111111111111001","000000000000000000","111111111111111011","111111111111110100","000000000000000000","111111111111011110","000000000000000000","111111111111100111","000000000000101110","000000000000010110","000000000000010101","111111111111111110","111111111111110101","111111111111111000","111111111111101111","111111111111110011","000000000000000011","000000000000000101","000000000000000101","000000000000010110","000000000000001001","000000000000000011","000000000000000000","111111111111110000","000000000000010111","111111111111111000","111111111111110110","111111111111111111","000000000000001000","000000000000000101","000000000000101111","111111111111010111","000000000000011001","111111111111111010","000000000000000010"),
("000000000000001001","000000000000000010","000000000000010110","111111111111100101","111111111111010011","000000000000000000","111111111111101101","111111111111111000","111111111111110100","000000000000101010","000000000000101100","000000000000011110","000000000000100000","111111111111110110","111111111111110110","111111111111101001","111111111111011111","111111111111111011","111111111111110101","111111111111100101","000000000000011111","000000000000000110","111111111111110010","000000000000001110","000000000000100100","000000000000001011","000000000000001111","111111111111110101","111111111111101110","111111111111100011","000000000000001111","111111111111110011","000000000000000000","000000000000011000","000000000000001001","111111111111110101","111111111111110011","111111111111110010","000000000000000101","111111111111111101","000000000000101110","111111111111111110","000000000000001010","111111111111110110","000000000000000111","000000000000000001","111111111111111111","000000000000001000","000000000000100001","111111111111011010","111111111111101110","000000000000000011","000000000000001010","000000000000010011","111111111111110100","000000000000100000","000000000000001010","000000000000000011","000000000000010101","111111111111111110","000000000000011011","111111111110001011","111111111110110100","000000000000000010","000000000000000111","111111111111111110","111111111111011000","000000000000000001","000000000000011010","000000000000011001","000000000000000111","000000000000000011","000000000000000101","000000000000000100","000000000000010000","111111111111100011","000000000000011100","111111111111110100","111111111111110111","111111111111101111","111111111111111100","000000000000000101","000000000000001100","111111111111110100","000000000000000101","111111111111111110","000000000000001101","111111111111111011","000000000000001100","111111111111101010","000000000000011100","111111111111111011","111111111111101011","000000000000000000","000000000000001110","000000000000000010","000000000000010100","000000000000000000","111111111111011001","000000000000001010","111111111111110110","000000000000001110","000000000000001101","000000000000000111","000000000000011011","111111111111110011","000000000000000101","111111111111110011","111111111111110001","000000000000000001","000000000000001111","111111111111111100","111111111111101100","000000000000001100","111111111111111111","000000000000000001","000000000000000101","000000000000001000","000000000000000010","000000000000000110","111111111111110000","000000000000101110","111111111111101010","000000000000010101","111111111111110100","000000000000000011","000000000000000010","000000000000010101"),
("000000000000100011","111111111111111101","000000000000100000","111111111111110001","111111111111001110","000000000000010010","111111111111101110","000000000000000001","111111111111110100","000000000000101011","000000000000101010","111111111111110011","111111111111110001","111111111111110001","111111111111110110","111111111111101010","111111111111100001","111111111111101000","000000000000000011","111111111111010111","000000000000100111","111111111111111010","111111111111110111","000000000000100011","000000000000001000","000000000000010001","000000000000001010","111111111111101111","111111111111001100","111111111111101011","111111111111111101","111111111111101100","000000000000001011","000000000000001110","000000000000010000","000000000000000000","111111111111111000","000000000000001111","000000000000011100","000000000000001110","000000000000010101","000000000000001011","111111111111101110","111111111111110001","000000000000100010","111111111111111100","111111111111100011","111111111111111111","000000000000000000","111111111111001101","111111111111110100","000000000000010010","000000000000000111","000000000000010110","111111111111111100","000000000000000000","000000000000010101","000000000000000000","000000000000001101","111111111111111001","000000000000001010","111111111110011111","111111111111000110","111111111111110001","000000000000001101","111111111111111000","000000000000100001","000000000000000110","111111111111110111","000000000000101111","000000000000010010","000000000000000100","111111111111111001","111111111111110110","111111111111110101","111111111111101000","000000000000001100","111111111111110011","000000000000001111","000000000000000011","000000000000011101","000000000000001110","000000000000001001","111111111110110000","000000000000001101","000000000000010001","000000000000011011","111111111111111011","111111111111110100","111111111111111100","000000000000011111","111111111111111001","111111111111111001","111111111111111000","111111111111101100","000000000000000101","000000000000010001","111111111111111100","111111111111111100","111111111111101011","111111111111111000","111111111111101011","000000000000011101","111111111111110111","000000000000101000","111111111111110110","000000000000001101","111111111111101000","111111111111101100","000000000000001111","000000000000011000","111111111111100101","111111111111110100","000000000000000010","111111111111101110","000000000000010001","111111111111101010","000000000000101010","000000000000011110","111111111111110011","111111111111110111","000000000000101101","111111111111111011","000000000000110110","111111111111111001","000000000000000101","111111111111110000","111111111111111100"),
("000000000000010110","111111111111011111","111111111111111000","111111111111011101","111111111111000000","111111111111110001","111111111111110011","000000000000001011","000000000000010111","000000000001000111","000000000000010010","000000000000000100","000000000000000101","000000000000010001","111111111111000101","111111111111111001","111111111111001011","111111111111011110","000000000000010010","111111111111110110","000000000001010011","111111111111100111","111111111111100010","000000000000100100","000000000000001000","111111111111111011","111111111111010111","111111111111110101","111111111111100111","000000000000010001","111111111111110000","000000000000010001","111111111111011111","000000000000010111","000000000000010111","111111111111011111","111111111111111111","000000000000001110","111111111111011111","000000000000010111","000000000000101110","000000000000100101","000000000000010100","000000000000011011","000000000000001001","000000000000010111","111111111111110001","111111111111011010","000000000000001000","111111111111101110","000000000000001100","111111111111111011","111111111111111110","000000000000010000","111111111111111100","000000000000001101","000000000000000110","000000000000010100","000000000000100011","111111111111101101","000000000000000110","111111111101110001","111111111111001110","111111111111011111","000000000000001001","111111111111111001","000000000000100011","000000000000001000","000000000000000110","000000000000001011","000000000000010110","000000000000000000","000000000000100011","000000000000011110","000000000000001010","111111111111110000","111111111111100011","111111111111101011","111111111111110001","111111111111111101","111111111111110110","111111111111110101","111111111111111000","111111111110001110","000000000000010001","000000000000111001","111111111111111101","111111111111111111","111111111111110000","000000000000100111","000000000000001111","111111111111111010","000000000000000010","000000000000010001","000000000000001000","111111111111111111","000000000000100010","111111111111110010","000000000000101111","111111111111100001","111111111111111011","111111111110011100","000000000000010001","111111111111101101","000000000000100000","111111111111110011","111111111111111010","111111111111101110","111111111111011111","111111111111100111","000000000000100011","111111111111101110","111111111111111011","000000000000010000","111111111111110001","111111111111101001","111111111111101100","000000000000100111","111111111111111110","000000000000000010","111111111111111011","000000000000010111","000000000000000101","000000000000100111","000000000000010111","111111111111100100","111111111111100110","111111111111110011"),
("111111111111101010","111111111111001111","111111111111110010","111111111111101111","000000000000000000","111111111111111101","111111111111111001","111111111111111100","000000000000011100","111111111111111101","000000000000000111","111111111111100110","000000000000001111","000000000000000101","111111111111010101","111111111111101101","111111111111001011","000000000000000110","000000000000011110","000000000000000111","000000000001010101","111111111111110110","111111111110111101","000000000000001010","111111111111111111","000000000000010000","111111111110111101","111111111111110111","111111111111111000","111111111111111101","111111111111110010","111111111111101000","000000000000000000","000000000000000000","000000000000101000","000000000000000001","000000000000001100","000000000000100010","111111111111010011","000000000000001111","000000000000010100","000000000000000100","000000000000001101","000000000000001001","111111111111101010","000000000000010101","000000000000000011","111111111110111011","111111111111101111","000000000000100001","000000000000010110","111111111111111010","111111111111111110","000000000000001011","000000000000000110","000000000000001000","111111111111011111","000000000000001000","000000000000011110","111111111111101101","000000000000010000","111111111110010101","111111111111100110","111111111111011100","000000000001001011","000000000000001001","000000000000100011","111111111111101101","111111111111111110","000000000000000000","111111111111111010","000000000000000000","000000000000101100","000000000000110011","000000000000010010","000000000000001001","111111111111111101","111111111111010100","000000000000001100","111111111111111111","111111111111111111","111111111111100110","111111111111010100","111111111111001101","000000000000001111","000000000000011010","111111111111100011","111111111111110111","000000000000000000","000000000000111001","111111111111111010","000000000000000000","000000000000101101","000000000000011111","111111111111111100","111111111111011000","000000000000110101","111111111111111001","000000000000111001","111111111111100000","111111111111111010","111111111110110010","000000000000000010","111111111111111110","000000000000110011","000000000000000001","000000000000011100","111111111111101000","111111111111000011","111111111111110111","000000000000011111","111111111111011001","111111111111101111","000000000000011011","111111111111100100","111111111111101111","111111111111110010","000000000000011000","111111111111110100","111111111111111110","111111111111011010","111111111111101111","000000000000010001","111111111111101001","000000000000000111","111111111111011101","111111111111101110","000000000000000111"),
("111111111111100010","111111111111101111","000000000000001000","111111111111110101","000000000001001111","111111111111111000","111111111111011000","111111111111111010","000000000000011111","111111111111011111","000000000000000101","111111111111101001","000000000000010000","000000000001001000","000000000000000100","111111111111101010","111111111111110010","111111111111100101","000000000000001101","000000000000000000","000000000000110100","000000000000000010","111111111111000011","000000000000011100","111111111111111000","000000000000001010","111111111111100101","111111111111101110","000000000000100100","000000000000000110","000000000000000001","000000000000000000","111111111111011110","111111111111100000","000000000000110000","000000000000010001","000000000000000001","000000000000001101","111111111111101110","000000000000000111","111111111111111011","000000000000010000","000000000000010110","000000000000011000","111111111111111010","000000000000101011","000000000000001101","111111111111010011","000000000000000011","111111111111111110","000000000000000100","111111111111111010","000000000000001001","000000000000001111","000000000000001110","111111111111111011","111111111111011100","000000000000001010","111111111111111111","111111111111101111","000000000000010110","111111111111110001","111111111111110000","111111111111111001","000000000000100011","111111111111110001","000000000000100101","111111111111010100","111111111111101001","111111111111011111","111111111111111011","000000000000001000","000000000000110011","000000000000110111","111111111111101100","111111111111111101","111111111111110110","111111111111101010","000000000000001000","111111111111101000","111111111111110100","111111111111110011","111111111111011110","000000000000011100","111111111111111001","000000000000011010","111111111111101010","111111111111111111","111111111111111111","000000000000101001","111111111111010011","111111111111110101","000000000000111110","000000000000011110","000000000000010011","111111111111010010","000000000000101010","000000000000000011","000000000000000110","111111111110110000","111111111111101011","111111111111100100","111111111111100010","000000000000001000","000000000000011011","000000000000001000","000000000000100101","111111111111011001","111111111111110011","111111111111101101","000000000000001011","111111111111111100","111111111111111101","000000000000000000","111111111111010001","111111111111101001","111111111111101101","000000000000011011","000000000000001000","111111111111111001","111111111111010010","111111111111101011","111111111111111101","111111111111100011","000000000000011110","111111111111000000","111111111111100011","000000000000000000"),
("111111111111000010","000000000000000111","000000000000010011","000000000000010001","000000000001000010","111111111111011111","111111111111100010","111111111111101010","000000000000010111","111111111111100101","111111111111100000","111111111111110011","000000000000001001","000000000000110001","111111111111110010","111111111111111110","000000000000011010","000000000000001010","000000000000000000","111111111111110011","000000000001000010","000000000000000011","000000000000010100","111111111111101101","000000000000010011","000000000000000100","000000000000001111","111111111111111100","000000000000101100","111111111111111011","111111111111101100","111111111111111101","111111111111111110","111111111111001100","000000000000000011","000000000000010110","111111111111101101","000000000000001011","111111111111101000","000000000000001111","111111111111011001","111111111111111011","000000000000010101","000000000000101001","111111111111100010","000000000000001100","111111111111110101","111111111111101000","000000000000001101","000000000000100101","111111111111110101","111111111111101001","111111111111110000","111111111111111100","000000000000001000","111111111111111000","111111111111101101","000000000000101000","000000000000000000","000000000000000101","000000000000011000","000000000000110001","000000000000001011","000000000000000111","000000000000010111","111111111111111011","000000000000000110","111111111111111000","111111111111111101","000000000000000011","000000000000000000","000000000000000101","000000000001001001","000000000000110010","111111111111101010","000000000000000100","000000000000000010","111111111111110001","111111111111110000","000000000000001111","111111111111101111","111111111111111010","111111111111111101","000000000000100001","111111111111111010","000000000000000000","111111111111110001","111111111111111011","111111111111100100","000000000000000101","111111111111010010","111111111111110110","000000000001001110","111111111111110100","000000000000010010","111111111111101100","000000000000010000","000000000000001011","111111111111111100","111111111110101010","111111111111101011","111111111111110000","111111111111111000","000000000000000010","000000000000001010","000000000000001111","000000000000000100","111111111111100100","000000000000101011","000000000000000010","111111111111111010","000000000000000110","111111111111011110","000000000000000000","111111111111111110","111111111111111011","111111111111101001","000000000000010001","000000000000000100","000000000000000110","111111111111001001","111111111111111000","111111111111110011","111111111111111100","000000000000011110","111111111111100100","111111111111011100","111111111111111011"),
("111111111110111001","000000000000001001","000000000000010010","111111111111111000","000000000000101110","111111111111110010","000000000000000000","000000000000000111","000000000000100010","111111111111111111","111111111111101111","111111111111101110","000000000000001110","000000000000010010","111111111111101110","111111111111110001","000000000000111110","000000000000000000","000000000000001010","000000000000010100","000000000000010100","000000000000000011","000000000000111001","000000000000000100","000000000000010010","000000000000000111","000000000000001101","000000000000000001","000000000000101110","111111111111100011","111111111111110010","000000000000010001","111111111111111000","111111111111000001","111111111111111011","000000000000011010","000000000000000000","000000000000001000","111111111111111001","000000000000001001","111111111111110010","111111111111011101","000000000000100001","000000000000011010","000000000000010100","111111111111111110","111111111111111001","111111111111101001","000000000000000011","000000000000001111","000000000000011110","000000000000001111","000000000000010100","111111111111101011","000000000000001000","111111111111111000","111111111111011011","000000000000100000","000000000000001010","000000000000001011","111111111111111111","000000000000101001","000000000000100010","000000000000000000","111111111111110110","111111111111101101","000000000000011100","111111111111101100","111111111111111001","000000000000101010","000000000000000000","111111111111110010","000000000000001011","000000000000110100","111111111111110011","111111111111110010","111111111111101011","111111111111111111","111111111111110111","000000000000001100","000000000000000110","000000000000001100","111111111111111101","000000000000100000","111111111111111000","000000000000010000","111111111111010011","111111111111100110","111111111111110101","111111111111101001","111111111111011100","111111111111110011","000000000001000110","111111111111110001","000000000000011010","111111111111110011","000000000000001001","111111111111100001","111111111111101101","000000000000000000","000000000000000011","111111111111011010","111111111111101010","111111111111110101","111111111111111010","000000000000000011","000000000000011011","111111111111111011","000000000000011101","000000000000001111","000000000000000000","000000000000000100","111111111111111100","111111111111111000","111111111111101111","111111111111010011","111111111111110010","000000000000010001","000000000000000000","000000000000000111","111111111111010110","111111111111101100","111111111111100100","111111111111111011","111111111111110100","111111111111110010","111111111111100001","000000000000010001"),
("111111111110110011","111111111111100011","000000000000010101","000000000000001100","111111111111100010","000000000000000010","111111111111111010","000000000000100100","000000000000000010","000000000000001111","000000000000010100","111111111111111001","111111111111111101","000000000000010011","000000000000001100","000000000000000111","000000000000100111","111111111111110010","111111111111111100","000000000000010001","000000000000001100","000000000000000011","000000000000111011","111111111111110101","000000000000010010","111111111111110100","000000000000001111","000000000000100011","000000000000011011","111111111111110001","000000000000000010","000000000000001001","000000000000010010","111111111111000011","111111111111101110","000000000000011101","111111111111100000","111111111111101111","000000000000001111","111111111111110010","111111111111111010","111111111111100000","111111111111110111","000000000000010011","000000000000000100","111111111111100111","000000000000000101","111111111111011010","000000000000010110","000000000000011100","000000000000000010","000000000000001010","000000000000000000","111111111111101100","000000000000000110","111111111111111111","111111111111110000","000000000000010010","000000000000100100","111111111111101101","111111111111111101","111111111111101110","000000000000000100","000000000000001000","111111111111110100","000000000000000000","000000000000010100","111111111111101110","111111111111101000","000000000000111101","000000000000000111","111111111111111011","000000000000001010","000000000000000100","000000000000000010","111111111111101011","111111111111111111","000000000000001000","000000000000001000","000000000000001110","111111111111111111","000000000000000010","000000000000000010","000000000000001100","000000000000001100","000000000000001001","111111111111100101","111111111111101001","111111111111100110","111111111111010010","111111111111100110","000000000000000100","000000000000111101","111111111111100011","000000000000100101","111111111111111110","111111111111011111","111111111111111010","000000000000000010","000000000000100001","111111111111111110","111111111111011100","111111111111111110","000000000000000011","000000000000100010","111111111111111010","000000000000011001","111111111111111001","000000000000001100","000000000000000110","000000000000001010","000000000000000111","000000000000001000","000000000000001101","000000000000000000","000000000000000000","000000000000001110","000000000000000000","000000000000010000","000000000000001110","111111111111010110","111111111111110100","111111111111111100","000000000000011101","000000000000001001","111111111111110110","111111111111100001","000000000000001011"),
("111111111111011001","111111111111101000","000000000000010000","000000000000001111","111111111111101111","000000000000010111","000000000000000000","000000000000010101","000000000000011001","111111111111111110","000000000000001000","111111111111101001","000000000000010101","000000000000100101","000000000000010001","000000000000000010","000000000000010110","111111111111110000","000000000000010010","000000000000001110","000000000000100101","000000000000001011","000000000000011010","000000000000001010","000000000000000100","111111111111110011","000000000000010010","000000000000011000","111111111111111010","111111111111011000","000000000000001100","000000000000001101","000000000000000000","111111111110110000","111111111111110000","000000000000100011","111111111111111111","000000000000010111","000000000000000110","000000000000001111","111111111111110000","111111111111110010","111111111111011100","000000000000010000","111111111111111010","111111111111101011","111111111111101000","111111111111111011","000000000000011010","000000000000001110","000000000000000100","111111111111111000","000000000000011110","111111111111100001","000000000000000000","000000000000001101","111111111111011001","000000000000010110","000000000000010111","111111111111101111","111111111111110001","111111111111111101","000000000000001001","000000000000100001","111111111111101011","111111111111101101","111111111111111000","111111111111110101","111111111111011110","000000000000011111","000000000000011000","111111111111110011","000000000000001101","000000000000000000","111111111111011100","111111111111111101","000000000000001011","000000000000010010","000000000000011011","000000000000000101","111111111111100101","000000000000001011","000000000000000111","000000000000001110","000000000000010100","000000000000010101","111111111111001101","111111111111100110","111111111111101000","111111111111001010","111111111111100010","111111111111101100","000000000001001011","111111111111101011","000000000000001100","111111111111111010","111111111110110001","111111111111110011","000000000000000011","000000000000111101","000000000000000101","000000000000000111","111111111111110101","000000000000100000","000000000000010100","000000000000100010","000000000000011111","111111111111111100","000000000000001111","111111111111101111","000000000000010101","000000000000000001","111111111111110100","111111111111111010","000000000000001100","000000000000000000","000000000000000100","000000000000010010","111111111111111001","111111111111101100","111111111110111010","111111111111111010","111111111111011100","000000000000000010","000000000000001101","111111111111111000","111111111111100110","000000000000010011"),
("111111111111011000","000000000000001000","111111111111111011","000000000000010001","111111111111001010","111111111111110001","000000000000010100","111111111111110101","111111111111111000","000000000000000001","000000000000100000","111111111111101100","111111111111101110","111111111111111101","000000000000000000","000000000000000000","111111111111100111","111111111111111110","111111111111110111","000000000000000101","000000000000010100","000000000000110000","000000000000010011","000000000000001001","111111111111111110","111111111111110001","000000000000100100","000000000000011001","111111111111100110","111111111111101101","111111111111111101","000000000000001101","000000000000000111","111111111111000100","000000000000000110","000000000000001011","111111111111110100","000000000000010101","000000000000001111","000000000000000000","111111111111101010","111111111111100001","111111111111001011","111111111111011000","111111111111110100","111111111111100110","111111111111110000","111111111111110001","000000000000100110","000000000000010011","111111111111111111","111111111111111010","000000000000100101","000000000000000000","111111111111101101","000000000000000100","111111111111100100","000000000000011000","000000000000001111","111111111111101101","000000000000010000","000000000000000011","000000000000011001","000000000000001001","111111111111001111","111111111111111011","000000000000011001","111111111111101100","111111111111111001","000000000000100101","111111111111111100","000000000000010110","000000000000101000","111111111111100000","111111111111011100","111111111111110011","111111111111111001","000000000000011100","000000000000000101","000000000000010001","111111111111110000","111111111111111010","000000000000010000","000000000000001110","111111111111111110","000000000000000101","111111111111110110","111111111111010101","111111111111011011","111111111111100110","111111111111101111","000000000000001111","000000000001001101","000000000000000010","111111111111111100","111111111111110111","111111111111011110","111111111111101101","111111111111111110","000000000001000001","000000000000000011","111111111111100110","000000000000001101","000000000000000111","000000000000010111","000000000000011101","000000000000010101","111111111111110101","000000000000000010","111111111111110111","000000000000000010","111111111111111011","111111111111101000","000000000000010100","000000000000110010","000000000000101001","000000000000000000","111111111111111111","111111111111111101","111111111111110010","111111111111001011","111111111111101011","111111111111100000","000000000000001111","111111111111101111","111111111111011111","111111111111110110","111111111111111000"),
("111111111111010010","111111111111011110","000000000000010011","000000000000001011","111111111111010010","000000000000000110","000000000000001111","111111111111011100","111111111111101011","000000000000011011","000000000000000000","000000000000000101","111111111111101011","000000000000000000","000000000000010011","111111111111110011","111111111111110111","000000000000000111","000000000000000010","111111111111111100","000000000000010001","000000000000101010","111111111111111010","000000000000001111","000000000000001010","111111111111101011","000000000000010101","111111111111111010","111111111111001100","000000000000001011","000000000000001010","111111111111111110","111111111111110100","111111111110011011","000000000000000111","111111111111101101","111111111111101011","111111111111101111","000000000000011100","000000000000001111","111111111111100011","111111111111011011","111111111111011111","111111111110111010","000000000000001000","111111111111111010","000000000000000011","111111111111100101","000000000000100100","000000000000000000","111111111111111101","000000000000000000","000000000000000111","111111111111011010","111111111111011110","000000000000100011","111111111111010110","000000000000000000","000000000000010110","111111111111110111","000000000000001110","111111111111101010","000000000000001110","111111111111111100","111111111111010101","000000000000000111","000000000000100100","111111111111101111","111111111111100001","000000000000010001","000000000000000000","000000000000101101","000000000000000001","111111111111010001","111111111111100111","111111111111100001","111111111111110010","000000000000011101","000000000000011101","000000000000100010","111111111111110010","111111111111110011","000000000000000011","111111111111110100","000000000000010000","111111111111110001","111111111111111101","111111111111011001","111111111111111110","111111111110111110","000000000000001010","111111111111111011","000000000000101110","000000000000001101","111111111111100001","111111111111101110","111111111111010101","000000000000001110","111111111111101110","000000000000111001","111111111111111000","111111111111110100","000000000000000100","000000000000010000","000000000000100010","000000000000001010","111111111111111010","111111111111110110","000000000000010011","000000000000000010","111111111111111101","000000000000011000","111111111111111001","000000000000000100","000000000000011101","000000000000010011","111111111111100111","000000000000010111","000000000000001001","000000000000010101","111111111111010101","000000000000011100","000000000000001001","000000000000011111","111111111111101111","111111111111010110","111111111111110100","000000000000000111"),
("111111111111001001","111111111111011111","000000000000000001","000000000000100000","111111111111110111","111111111111111001","000000000000001010","111111111111101011","111111111111110010","000000000000011101","111111111111110001","111111111111011101","000000000000000100","111111111111110100","000000000000001111","000000000000000001","111111111111110000","000000000000001110","000000000000001100","000000000000011100","000000000000100001","000000000000111011","111111111111111111","000000000000001010","111111111111111010","111111111111111010","000000000000000000","111111111111111001","111111111111101011","000000000000001010","111111111111111100","000000000000100010","000000000000001101","111111111110101101","111111111111101110","111111111111011000","111111111111101111","111111111111110001","000000000000100000","111111111111110101","111111111111111011","111111111111111010","111111111111101101","111111111111010011","111111111111110110","111111111111101000","000000000000000110","111111111111100010","000000000000011010","000000000000001101","000000000000101100","000000000000000101","000000000000011001","111111111111111100","111111111111111001","000000000000010011","111111111111100001","000000000000011000","000000000000001100","111111111111111011","000000000000011011","111111111111110111","111111111111101001","111111111111110001","111111111111101010","000000000000001011","000000000000110001","111111111111011101","111111111111100011","111111111111110110","111111111111101100","000000000000011010","000000000000101001","111111111110111110","111111111111100110","111111111111111111","111111111111100001","000000000000001001","000000000000000100","000000000000101110","000000000000001101","111111111111111101","000000000000000100","111111111111111001","000000000000010011","111111111111100011","111111111111110101","111111111110111001","111111111111011100","111111111111101101","111111111111111110","000000000000000001","000000000000001101","000000000000001001","111111111111100100","111111111111111110","111111111111011011","111111111111111010","000000000000001000","000000000000011100","111111111111011110","000000000000000001","000000000000010010","000000000000000000","111111111111111101","000000000000100111","111111111111111111","000000000000000101","000000000000000111","111111111111110010","000000000000001101","000000000000010011","000000000000000000","000000000000010000","000000000000110001","000000000000100110","000000000000000001","000000000000010100","000000000000010000","000000000000010001","111111111111011000","111111111111101110","000000000000000010","000000000000011110","111111111111111001","111111111111001011","111111111111111010","000000000000000010"),
("111111111111100110","000000000000000011","111111111111101000","000000000000000101","111111111111111001","111111111111100010","000000000000000001","000000000000000111","000000000000001110","000000000000101000","000000000000001110","111111111111111100","111111111111100111","111111111111111100","111111111111111000","000000000000001011","111111111111001101","000000000000001111","000000000000000100","111111111111111011","000000000000001010","000000000000010010","000000000000000000","000000000000011010","111111111111111101","000000000000001111","000000000000100010","000000000000000011","111111111111100000","000000000000000101","111111111111111011","000000000000000000","000000000000001100","111111111111100000","111111111111110110","111111111111101101","111111111111100100","111111111111101001","000000000000011000","111111111111101100","111111111111110010","000000000000000110","111111111111100100","111111111111001100","000000000000000100","111111111111110000","111111111111111000","111111111111101010","111111111111111011","111111111111110010","000000000000010011","000000000000011111","000000000000010010","111111111111101110","111111111111110111","000000000000000101","000000000000001101","000000000000001110","000000000000010001","000000000000001111","000000000000011110","000000000000000001","111111111111010011","000000000000000111","111111111111010110","111111111111101001","000000000000101000","111111111111111001","111111111111111110","111111111111111101","000000000000000101","111111111111111100","000000000000110111","111111111110111000","000000000000000000","000000000000000001","111111111111110101","111111111111110000","111111111111111100","000000000000001010","000000000000000001","000000000000000010","111111111111110110","111111111111001110","000000000000011101","111111111111111000","111111111111101000","111111111111100000","111111111111110110","111111111111100101","111111111111100001","000000000000101001","000000000000010111","000000000000010100","111111111111101010","000000000000000111","111111111111110101","000000000000010001","000000000000011111","000000000000000101","111111111111100111","111111111111111110","000000000000101110","000000000000011011","000000000000010101","000000000000101011","000000000000001100","000000000000001110","111111111111111000","111111111111011100","000000000000011001","000000000000000100","000000000000001011","111111111111111101","000000000000001011","000000000000011001","000000000000001110","000000000000001101","000000000000011111","111111111111110001","111111111110111001","111111111111111110","111111111111010110","000000000000001110","111111111111100001","111111111111010111","111111111111101111","000000000000001110"),
("111111111111010000","000000000000000110","000000000000001011","111111111111011111","111111111110111011","111111111111111001","111111111111111101","111111111111110101","111111111111100101","000000000000000000","111111111111110101","000000000000000000","000000000000010010","000000000000010001","111111111111110010","000000000000000000","111111111111010010","000000000000000010","111111111111111100","111111111111111001","000000000000110111","111111111111111111","000000000000000000","000000000000000111","000000000000101000","111111111111110110","000000000000100001","111111111111010110","111111111111100010","000000000000101001","000000000000000000","111111111111100011","000000000000010011","111111111111011011","000000000000001110","111111111111011110","000000000000010100","111111111111110011","000000000000101111","111111111111111101","000000000000001110","000000000000001110","111111111111011010","111111111111010101","000000000000000011","111111111111110000","000000000000000111","000000000000010110","000000000000100000","111111111111010001","111111111111101111","000000000000101010","000000000000011110","111111111111100010","111111111111111011","111111111111110010","000000000000010100","111111111111010101","111111111111100111","000000000000000000","000000000000000111","111111111111101111","111111111110110111","111111111111100111","111111111111111001","000000000000110111","000000000000110101","000000000000001010","111111111111100110","000000000000001010","111111111111101101","111111111111111010","000000000000011111","111111111111000101","111111111111110011","111111111111101101","000000000000110000","111111111111100110","111111111111110100","111111111111110011","000000000000010000","000000000000001001","111111111111011011","111111111111011111","111111111111111011","111111111111111011","111111111111100010","111111111111111110","111111111111110010","111111111111010011","111111111111110000","000000000000010010","000000000001010011","000000000000000010","111111111111100001","111111111111110111","111111111111111100","000000000000001011","000000000000100110","111111111111111000","111111111111111101","000000000000000111","111111111111011111","111111111111111111","000000000000110001","000000000000000111","111111111111101101","000000000000011001","111111111111110000","111111111111110110","000000000000001101","000000000000000011","000000000000010000","111111111111001111","111111111111111100","111111111111101110","111111111111100110","111111111111110110","000000000001001010","111111111111101110","111111111111001110","000000000000010110","111111111111111011","000000000000001100","111111111111010101","111111111111111111","000000000000000110","111111111111111100"),
("000000000000010000","000000000000001111","000000000000101011","000000000000000011","111111111111001101","111111111111001111","111111111111111001","111111111111111100","111111111111111101","111111111111100101","111111111111111000","111111111111111001","000000000000011001","000000000000011111","111111111111111101","111111111111111010","111111111111101000","000000000000001101","000000000000000100","000000000000011001","000000000000010101","111111111111100111","111111111111101111","111111111111110111","000000000000001001","111111111111100110","000000000000100001","111111111111011001","111111111111101000","000000000000010110","000000000000011110","000000000000000100","000000000000000110","000000000000000010","000000000000001000","111111111111011110","000000000000000110","000000000000000101","000000000000100101","000000000000000011","000000000000000110","000000000000010011","111111111111111010","111111111111110011","000000000000010111","000000000000000000","111111111111101101","111111111111111101","000000000000101100","111111111111011010","111111111111110000","000000000000001111","111111111111111001","000000000000000000","000000000000000000","111111111111110100","000000000000101101","111111111111110011","111111111111011100","111111111111110110","000000000000000110","000000000000010011","111111111111110001","111111111111101011","111111111111101000","000000000000011101","000000000000101011","111111111111011111","000000000000000011","000000000000010011","111111111111010010","111111111111111101","000000000000110000","111111111111111101","111111111111101101","000000000000010010","000000000000001110","111111111111100110","111111111111101010","111111111111100011","000000000000011000","000000000000100011","111111111111011110","111111111111101111","000000000000001100","111111111111100111","000000000000010100","000000000000010001","111111111111101011","000000000000000110","111111111111111111","111111111111100100","000000000000101011","111111111111000001","111111111111101110","111111111111100110","000000000000100010","000000000000000000","000000000000001101","111111111111111111","000000000000010000","111111111111101001","111111111111010010","111111111111100111","000000000000010111","111111111111011111","000000000000000000","000000000000001100","000000000000001011","111111111111110101","000000000000010001","000000000000000010","111111111111101001","111111111111101110","000000000000000010","111111111111000011","111111111111010101","000000000000000100","000000000000110101","000000000000001111","111111111111111011","000000000000001100","000000000000000000","111111111111011000","111111111111011100","111111111111111100","000000000000100011","000000000000110011"),
("111111111111110111","111111111111011011","000000000000011101","000000000000001010","111111111111101100","111111111111111101","111111111111101001","111111111111100110","000000000000000111","111111111111001010","000000000000000000","000000000000010110","000000000000001010","111111111111110010","111111111111101011","111111111111111100","111111111111010100","000000000000001101","000000000000011001","000000000000000000","000000000000101100","111111111111011100","111111111111011110","111111111111100000","000000000000010010","000000000000000000","000000000000011010","111111111111100110","111111111111111100","000000000000001101","000000000000010011","111111111111111010","000000000000010000","000000000000000111","000000000000110110","111111111111100111","000000000000000110","000000000000011001","000000000000001101","000000000000001001","000000000000011011","000000000000101000","000000000000011100","000000000000000110","000000000000010001","111111111111100011","000000000000000000","000000000000001000","000000000000100111","111111111111110101","000000000000000101","000000000000101001","000000000000000110","000000000000100101","000000000000000000","111111111111111010","000000000000001010","111111111111100110","111111111111010110","111111111111101101","000000000000010111","000000000000000000","000000000000000101","111111111111100010","000000000000010000","000000000000010000","000000000000011111","111111111111111101","000000000000011100","000000000000100110","111111111111101010","000000000000001100","000000000000100101","111111111111110000","111111111111101101","000000000000001100","000000000000001000","111111111111110101","111111111111100101","111111111111100010","111111111111111010","111111111111111000","111111111111100011","111111111111110011","000000000000001110","111111111111111010","000000000000100000","111111111111111001","111111111111001111","000000000000010000","111111111111100110","111111111111110110","000000000000101000","111111111111101111","111111111111111100","111111111111010110","000000000000000111","000000000000011011","000000000000010001","111111111111110001","000000000000010110","111111111111101110","111111111111111000","111111111111111111","000000000000011101","111111111111101001","111111111111110110","111111111111110001","111111111111101010","111111111111011110","000000000000001001","000000000000000000","000000000000000011","000000000000010001","111111111111111101","111111111111101011","111111111111011101","000000000000001011","111111111111111100","000000000000010111","000000000000000110","000000000000001011","000000000000000000","111111111111101010","111111111111110101","000000000000010110","000000000000101110","000000000000011001"),
("111111111111111001","000000000000010101","111111111111111110","111111111111110011","000000000000011100","111111111111101110","000000000000000001","111111111111111011","000000000000010001","111111111111101000","000000000000000011","000000000000000100","000000000000100100","000000000000010011","000000000000000000","000000000000001000","111111111111110101","000000000000000111","000000000000001001","111111111111110100","000000000000100000","000000000000001011","000000000000001110","000000000000010011","111111111111110011","111111111111111001","000000000000000001","111111111111110011","111111111111111011","111111111111101101","111111111111111001","000000000000001100","111111111111110001","000000000000000010","111111111111111001","000000000000001001","000000000000010000","111111111111100111","111111111111011001","000000000000011001","000000000000010101","000000000000010100","000000000000010011","111111111111111010","111111111111011011","000000000000000111","000000000000100010","111111111111111011","000000000000100001","000000000000001010","111111111111111110","111111111111111101","000000000000010001","000000000000001111","111111111111101101","000000000000001001","111111111111111101","111111111111101110","000000000000101001","000000000000010000","111111111111100011","000000000000010101","000000000000001010","111111111111100011","000000000000011000","000000000000010110","111111111111100011","111111111111011000","000000000000110110","111111111111111101","111111111111110111","000000000000001010","000000000000001010","111111111111110110","111111111111110101","111111111111111101","000000000000000001","000000000000000000","000000000000010010","000000000000010010","111111111111001111","111111111111011111","111111111111100101","000000000000010011","000000000000000100","000000000000010110","000000000000010000","111111111111111010","111111111111010111","000000000000010000","111111111111111101","111111111111110110","111111111111011111","111111111111111000","000000000000011000","000000000000000101","111111111111111111","111111111111100011","000000000000000000","000000000000111001","111111111111100111","111111111111101001","111111111111110110","000000000000000010","000000000000000000","000000000000000111","000000000000001000","000000000000000111","000000000000010000","111111111111101001","000000000000010100","111111111111110101","000000000000000010","111111111111111110","000000000000001101","000000000000001101","111111111111101011","000000000000000000","000000000000000011","000000000000010111","111111111111110110","111111111111101001","000000000000011111","111111111111111101","111111111111111000","111111111111100010","000000000000011010","000000000000011011"),
("111111111111110011","000000000000011000","000000000000001110","000000000000000011","111111111111110111","111111111111100110","000000000000001111","111111111111101001","000000000000000011","000000000000001111","111111111111011011","000000000000001001","000000000000000011","000000000000010110","000000000000001010","000000000000000001","000000000000001100","111111111111110110","000000000000000000","000000000000000010","000000000000010011","000000000000001000","000000000000000000","000000000000000111","000000000000101000","111111111111101110","000000000000001010","111111111111101100","000000000000000011","000000000000000100","111111111111111100","000000000000010100","111111111111110011","000000000000000010","000000000000010110","111111111111110001","000000000000001100","111111111111101100","111111111111111010","000000000000100101","000000000000011010","000000000000010101","000000000000000110","111111111111101001","111111111111011110","000000000000000000","000000000000011001","111111111111101100","000000000000010011","000000000000010111","111111111111111010","111111111111111000","111111111111111011","000000000000000101","111111111111111100","000000000000010001","000000000000000010","000000000000001001","000000000000010000","111111111111111100","111111111111111011","111111111111101110","111111111111111101","111111111111101111","111111111111100110","000000000000001001","111111111111110111","111111111111110111","000000000000011100","000000000000100010","111111111111111010","000000000000001000","000000000000001011","000000000000001001","111111111111110000","111111111111111100","111111111111110010","111111111111100001","000000000000100000","111111111111111000","000000000000000110","111111111111110100","111111111111111000","000000000000000110","111111111111111001","000000000000000010","000000000000100100","111111111111111011","000000000000000000","000000000000001001","000000000000000000","111111111111100111","000000000000010100","000000000000000010","000000000000000100","000000000000000000","000000000000001001","111111111111101010","000000000000001110","000000000000010011","000000000000001101","111111111111101010","000000000000001011","111111111111010111","111111111111111001","111111111111110110","000000000000010000","000000000000101001","000000000000001101","000000000000100001","000000000000011100","111111111111101101","111111111111101001","000000000000011000","000000000000000011","000000000000000101","111111111111100000","000000000000010000","111111111111110100","111111111111101100","000000000000011010","111111111111101100","111111111111110001","000000000000001110","000000000000011011","000000000000001000","000000000000001000","111111111111111011"),
("111111111111011100","000000000000000011","111111111111110111","111111111111101111","000000000000000100","111111111111101101","111111111111110010","111111111111010110","111111111111101000","000000000000100000","000000000000000111","111111111111111010","000000000000000000","000000000000000010","111111111111111010","111111111111110000","000000000000010000","000000000000001101","000000000000011010","000000000000011110","000000000000001011","000000000000011100","000000000000110000","000000000000100001","000000000000000101","111111111111100110","000000000000010111","111111111111101011","000000000000000111","111111111111111001","111111111111110101","000000000000011011","000000000000000001","000000000000001010","000000000000001011","111111111111100110","111111111111111101","000000000000001000","111111111111101111","000000000000001000","000000000000000101","000000000000000001","000000000000010101","000000000000011001","111111111111100010","000000000000010011","000000000000001111","000000000000010001","111111111111111110","000000000000000011","000000000000010100","000000000000010000","000000000000100011","000000000000001100","111111111111110110","111111111111011011","111111111111100101","000000000000000101","000000000000011101","111111111111110101","000000000000010101","000000000000000111","000000000000100100","111111111111101111","111111111111111101","000000000000011000","000000000000010111","111111111111111100","000000000000110100","000000000000101000","111111111111101001","000000000000001100","111111111111111011","000000000000000011","111111111111111111","000000000000000011","111111111111110001","111111111111111101","000000000000000010","000000000000001001","000000000000001001","111111111111101011","111111111111101000","000000000000001110","111111111111100100","000000000000010011","000000000000010110","000000000000000111","111111111111100101","000000000000010101","111111111111111000","111111111111111101","000000000000010100","000000000000100100","111111111111111111","000000000000000000","111111111111100011","111111111111010001","111111111111111000","111111111111110100","000000000000000010","111111111111110110","111111111111111111","111111111111111111","111111111111111111","000000000000101101","111111111111101000","111111111111111001","111111111111110110","000000000000011110","111111111111110100","111111111111101000","111111111111101001","000000000000001111","111111111111011101","000000000000011000","111111111111100100","000000000000011111","111111111111110011","000000000000001011","000000000000010011","000000000000010010","111111111111101000","000000000000000111","000000000000011001","111111111111101010","000000000000001100","111111111111010000"),
("000000000000000110","111111111111101111","000000000000001000","111111111111111001","000000000000001001","111111111111100011","111111111111101110","111111111111010010","000000000000010100","000000000000011100","111111111111100010","111111111111110110","000000000000000110","000000000000001111","000000000000101000","111111111111101100","000000000000001101","111111111111111111","000000000000010100","111111111111111010","000000000000100010","000000000000100010","111111111111110100","111111111111100100","000000000000010111","111111111111101111","111111111111101011","111111111111111100","000000000000011010","000000000000010101","111111111111011000","000000000000011110","111111111111101011","000000000000000111","000000000000000101","111111111111011111","111111111111111111","000000000000000111","111111111111100100","000000000000101111","000000000000010011","000000000000000110","000000000000001101","111111111111010011","111111111111111011","111111111111110001","111111111111111101","111111111111100010","000000000000100111","000000000000010001","111111111111111101","000000000000000100","000000000000100010","111111111111110000","111111111111111000","000000000000010100","111111111111111000","000000000000011100","000000000000000010","000000000000001111","000000000000001101","111111111111101011","111111111111010000","111111111111101101","000000000000001100","000000000000011111","000000000000010001","111111111111111001","111111111111111011","000000000000010000","111111111111101000","111111111111111101","000000000000000010","000000000000001100","111111111111101011","111111111111011111","111111111111100010","111111111111110000","000000000000100001","000000000000011011","111111111111011110","111111111111110011","111111111111110001","000000000000011111","111111111111100010","000000000000001011","000000000000100010","000000000000000011","111111111111110000","000000000000001010","111111111111111000","111111111111110010","000000000000011000","111111111111110101","000000000000011011","000000000000000110","111111111111111101","111111111111111010","000000000000000100","000000000000001101","111111111111111001","111111111111100011","000000000000001010","111111111111011010","000000000000000000","111111111111110010","111111111111111100","000000000000011000","111111111111110101","000000000000001010","000000000000011010","111111111111110101","111111111111110001","000000000000100000","000000000000011001","000000000000010000","111111111111111111","111111111111111100","111111111111011111","000000000000010001","000000000000001010","111111111111111011","000000000000000111","000000000000011011","000000000000010100","111111111111011010","000000000000000000","111111111111100011"),
("111111111111110100","111111111111110010","111111111111110111","111111111111111000","000000000000000001","111111111111101100","000000000000001011","000000000000101111","000000000000100101","000000000000001000","000000000000000100","000000000000000110","000000000000000111","111111111111111001","000000000000000000","111111111111110011","000000000000000000","000000000000010001","111111111111111100","000000000000011110","000000000000000101","111111111111111101","111111111111110000","111111111111111110","111111111111110111","000000000000000000","111111111111101101","000000000000001001","000000000000001001","111111111111111110","111111111111011111","000000000000101110","000000000000000001","000000000000000100","111111111111111101","111111111111110111","000000000000000001","000000000000000101","111111111111111011","000000000000000010","000000000000001011","111111111111101001","000000000000100101","111111111111110100","111111111111111000","000000000000000100","000000000000001001","111111111111100011","000000000000100010","000000000000101111","000000000000000101","111111111111101100","000000000000001111","111111111111111100","000000000000001001","000000000000000000","111111111111011100","000000000000001101","111111111111111100","111111111111110100","000000000000001011","111111111111101100","111111111111011001","111111111111111100","111111111111100111","111111111111111111","000000000000010001","111111111111110100","111111111111111001","000000000000010010","000000000000100000","000000000000100111","111111111111111011","000000000000010110","000000000000000001","111111111111011001","111111111111100011","111111111111011111","111111111111101001","000000000000010111","111111111111101000","111111111111110010","111111111111110001","000000000000001000","000000000000001101","111111111111111110","111111111111101101","111111111111111100","111111111111101000","000000000000101110","111111111111110011","111111111111101111","000000000000000000","000000000000010111","000000000000001011","111111111111011111","111111111111111011","000000000000011000","000000000000101011","000000000000001100","000000000000000111","111111111111100101","111111111111100000","111111111111111100","111111111111101110","000000000000100101","000000000000000100","111111111111111010","111111111111101101","111111111111111110","000000000000001000","000000000000001100","000000000000000010","000000000000111100","000000000000010000","111111111111101110","000000000000000000","000000000000000111","111111111111001010","000000000000001110","111111111111101101","111111111111100101","111111111111011101","000000000000010001","000000000000000010","111111111111110101","111111111111101111","111111111111110100"),
("111111111111110011","111111111111110010","111111111111100001","111111111111110001","111111111111100100","000000000000000010","111111111111111010","000000000000100001","000000000000010000","111111111111101010","000000000000110101","000000000000010000","111111111111111110","111111111111110011","111111111111111010","111111111111100011","111111111111101010","000000000000001001","000000000000010011","111111111111101010","000000000000010000","000000000000010001","111111111111100111","111111111111110111","111111111111111011","111111111111111001","111111111111111000","111111111111111000","000000000000000000","111111111111101111","111111111111101110","000000000000011111","111111111111111001","111111111111101100","000000000000001100","000000000000001010","111111111111101000","000000000000010110","111111111111011011","111111111111101011","000000000000100101","000000000000001010","000000000000011111","111111111111111101","111111111111111110","111111111111101111","000000000000011001","111111111111100100","000000000000000111","000000000000001011","111111111111001011","111111111111100101","000000000000010110","000000000000101010","000000000000000111","000000000000001010","111111111111111111","111111111111111110","000000000000001011","111111111111110100","000000000000000001","111111111110110110","111111111111100011","111111111111100000","111111111111100110","111111111111110000","000000000000001001","111111111111110100","111111111111100100","111111111111110101","000000000000000000","000000000000001100","111111111111111111","000000000000010011","000000000000111000","111111111111100110","111111111111110100","000000000000001100","000000000000000110","111111111111011011","111111111111010111","111111111111101101","111111111111100101","111111111111110100","000000000000011101","111111111111100000","000000000000001110","000000000000000010","111111111111001110","111111111111100011","111111111111010111","111111111111101001","000000000000001111","111111111111110101","111111111111110011","111111111111010111","111111111111000101","000000000000010101","000000000000001000","000000000000100100","111111111111101011","111111111111101100","111111111111110111","000000000000100011","000000000000001010","111111111111111101","000000000000001101","000000000000001100","111111111111101100","111111111111110000","111111111111111111","000000000000001010","000000000000001111","000000000000100010","000000000000100011","000000000000000001","000000000000010001","000000000000000101","111111111111000101","111111111111111111","000000000000011111","111111111111100110","111111111111111011","000000000000100111","111111111111011110","111111111111010001","111111111111001111","111111111111110101"),
("000000000000000000","000000000000001111","000000000000001101","000000000000000011","111111111111101110","111111111111110100","000000000000001001","000000000000110000","111111111111101001","111111111111010011","000000000000110111","000000000000010001","000000000000011011","111111111111011100","000000000000010000","111111111111011011","111111111111110111","000000000000000000","111111111111101010","111111111111111100","111111111111111001","000000000000011100","111111111111101101","111111111111011101","000000000000000101","000000000000000110","000000000000010101","111111111111101110","111111111111111001","111111111111110001","000000000000010001","111111111111111011","000000000000001111","111111111111011010","111111111111100101","000000000000000110","000000000000000101","111111111111110100","000000000000000000","111111111111111001","000000000000001110","111111111111111000","000000000000011001","000000000000000000","111111111111111100","111111111111010100","000000000000010001","111111111111110011","000000000000000110","000000000000001011","111111111111000110","111111111111110000","000000000000001100","000000000000010110","000000000000000001","000000000000100111","111111111111100100","111111111111001011","111111111111110000","111111111111110010","111111111111111100","111111111111001000","111111111111010110","111111111111111100","111111111111100011","000000000000000100","111111111111100111","111111111111110110","000000000000010010","111111111111100010","000000000000000111","111111111111110011","111111111111111001","111111111111111101","000000000000011000","111111111111110100","000000000000001011","111111111111111110","000000000000010010","111111111111100110","000000000000000110","000000000000101011","111111111111111101","111111111111100111","111111111111111000","111111111111011101","000000000000001011","111111111111110001","111111111111010001","111111111111011101","111111111111100011","111111111111100101","000000000000000110","111111111111010001","000000000000011010","111111111111100110","111111111111110110","000000000000110100","111111111111100101","000000000000011101","000000000000001101","111111111111111110","111111111111011001","000000000000001100","111111111111111111","000000000000000010","000000000000011100","111111111111111101","111111111111101100","111111111111101010","000000000000101001","000000000000010110","000000000000001101","000000000000000000","000000000000010101","111111111111101100","000000000000000010","000000000000000101","111111111111010111","111111111111101001","000000000000011111","000000000000000000","000000000000000000","000000000000111010","111111111111100110","111111111111110101","111111111111110000","000000000000010110"),
("111111111111010100","000000000000010101","000000000000001011","111111111111110111","111111111111101111","111111111111110101","000000000000001011","111111111111101001","111111111111101100","111111111111101010","000000000000110010","000000000000101101","000000000000000001","111111111111110100","111111111111110011","000000000000000110","111111111111001100","000000000000000000","000000000000001101","111111111111110000","111111111111111100","000000000000100110","000000000000010011","111111111111010001","000000000000001110","111111111111110100","000000000000000011","111111111111110001","111111111111111010","111111111111101111","000000000000000000","111111111111111101","111111111111111111","111111111111101001","000000000000010001","111111111111110011","000000000000010100","111111111111101000","111111111111111100","111111111111110110","000000000000000011","111111111111101101","000000000000010100","000000000000001001","111111111111111111","111111111111011110","000000000000011101","111111111111011110","111111111111110001","111111111111101110","111111111111010010","111111111111111000","000000000000001110","000000000000010111","000000000000000000","000000000000011101","111111111111100010","111111111111110100","000000000000001001","111111111111101110","111111111111100101","111111111111000100","111111111111000111","000000000000011100","111111111111000000","000000000000011100","111111111111100100","000000000000100111","000000000000000110","111111111111110000","000000000000000000","111111111111010101","111111111111010001","111111111111111100","000000000000001101","000000000000000011","000000000000001011","000000000000001000","111111111111101111","111111111111111011","000000000000001000","000000000000010110","111111111111110110","111111111111100101","111111111111100011","111111111111011010","000000000000010110","111111111111010010","111111111111101100","111111111111010000","111111111111001100","000000000000000101","000000000000000000","111111111111100001","000000000000101010","111111111111101101","111111111111111011","000000000000001111","111111111111011001","000000000000100001","000000000000001101","000000000000010010","111111111111111100","000000000000010100","111111111111101110","000000000000000000","000000000000010011","111111111111110010","111111111111111110","000000000000000101","000000000000000110","000000000000100011","111111111111111111","111111111111101101","000000000000001011","111111111111111011","000000000000010111","000000000000010101","111111111111110000","111111111111110000","000000000000010001","000000000000000010","000000000000010011","000000000000011011","111111111111101110","000000000000100000","000000000000001010","000000000000010010"),
("111111111111100100","000000000000011001","000000000000010000","000000000000001101","111111111111111101","000000000000010011","000000000000010010","111111111111010100","111111111111100111","111111111111111110","000000000000111111","000000000000000000","111111111111111100","111111111111101010","111111111111111111","111111111111110000","111111111111110000","000000000000000110","000000000000010010","111111111111001011","000000000000010101","000000000000000001","000000000000001001","111111111111011000","000000000000001111","111111111111111011","000000000000000110","111111111111100001","111111111111111000","111111111111111001","111111111111110010","000000000000001011","111111111111101010","111111111111100110","000000000000001110","111111111111111010","111111111111111001","111111111111100010","000000000000000010","000000000000000001","000000000000100000","000000000000000001","111111111111111101","111111111111110001","111111111111110001","111111111111111100","000000000000011010","111111111111110110","000000000000000110","111111111111111100","111111111111101011","111111111111110100","000000000000101110","000000000000010111","111111111111011111","000000000000010100","000000000000000001","111111111111111100","000000000000010100","111111111111110010","111111111111111101","111111111110010110","111111111111000010","000000000000010000","111111111111101011","000000000000001011","111111111111100010","000000000000000001","111111111111111001","000000000000000100","000000000000001000","111111111111111000","111111111111110101","000000000000000101","000000000000000011","111111111111111111","000000000000010010","000000000000001011","000000000000010101","111111111111110100","111111111111111010","000000000000000001","111111111111110011","111111111111101110","111111111111100011","111111111111101101","000000000000011101","111111111111100110","000000000000000000","111111111111011101","111111111111011101","000000000000011011","000000000000000000","111111111111110101","000000000000101111","111111111111110011","000000000000001011","000000000000001011","111111111111111001","000000000000110000","000000000000000111","000000000000001101","111111111111110000","111111111111111110","111111111111100010","000000000000011100","000000000000011101","000000000000011100","111111111111101001","111111111111101101","000000000000001101","111111111111111100","111111111111101011","000000000000001000","111111111111110010","111111111111110010","000000000000000010","000000000000011010","000000000000000100","111111111111101100","111111111111111001","000000000000000111","000000000000001001","000000000000101101","111111111111110100","000000000000101011","000000000000000110","111111111111111100"),
("000000000000000000","000000000000010001","000000000000010101","000000000000001010","000000000000010011","111111111111101001","000000000000001111","111111111111110111","111111111111100011","111111111111111111","000000000000100100","000000000000001101","111111111111101011","000000000000010110","000000000000011101","111111111111100000","111111111111101000","000000000000000000","000000000000001001","111111111111101100","000000000000011001","000000000000011001","000000000000000000","111111111111011111","000000000000000101","111111111111110010","000000000000000001","111111111111110111","111111111111110001","111111111111110100","111111111111110111","000000000000001000","000000000000000110","111111111111110101","000000000000000110","111111111111101111","000000000000000100","111111111111110101","111111111111111110","111111111111101011","000000000000011101","000000000000010001","111111111111110011","111111111111110000","000000000000011010","111111111111011101","000000000000010010","111111111111101111","111111111111111111","000000000000010100","111111111111110011","111111111111110111","000000000000001011","000000000000010010","111111111111111011","000000000000011001","000000000000001001","111111111111110101","000000000000011011","111111111111101010","000000000000001101","111111111110011100","111111111111000000","000000000000011101","000000000000001000","000000000000011010","111111111111011001","000000000000010110","111111111111100010","111111111111111101","111111111111101111","111111111111110111","000000000000000000","111111111111110100","111111111111110110","000000000000000111","000000000000011010","111111111111111011","000000000000001010","111111111111100100","000000000000001001","000000000000011011","111111111111111110","000000000000000010","111111111111101010","111111111111111010","000000000000010001","111111111111101000","000000000000010101","111111111111010001","111111111111011011","000000000000011111","000000000000101110","111111111111110001","000000000000100011","000000000000100011","111111111111111011","000000000000101100","111111111111100110","000000000000101001","000000000000000111","000000000000101011","000000000000011000","111111111111110010","111111111111101000","111111111111110111","000000000000010111","111111111111111110","000000000000001100","000000000000000111","000000000000001101","000000000000000001","000000000000001100","111111111111100111","000000000000011010","000000000000011011","111111111111111011","000000000000010100","000000000000001111","111111111111100001","000000000000000101","111111111111110110","000000000000000001","000000000000101011","111111111111100101","000000000000001100","111111111111111010","111111111111111111"),
("000000000000000000","000000000000110111","000000000000010101","111111111111110110","000000000000010111","000000000000001010","000000000000001010","111111111111110010","111111111111100001","000000000000011000","000000000000011101","000000000000011010","111111111111101101","000000000000000001","000000000000000010","111111111111010010","111111111111101000","111111111111100101","000000000000000111","111111111111100001","000000000000001101","000000000000010110","000000000000000101","111111111111011100","000000000000001111","000000000000001011","000000000000001101","111111111111111111","111111111111100110","111111111111001100","111111111111111111","000000000000000001","111111111111101010","000000000000000010","000000000000001001","111111111111101011","111111111111111001","111111111111111001","111111111111110110","000000000000000111","000000000000001011","000000000000001101","111111111111110111","111111111111101101","000000000000001010","111111111111110111","000000000000011011","000000000000001000","000000000000001101","000000000000010001","111111111111110000","000000000000001101","000000000000011101","111111111111101110","111111111111110111","000000000000001100","000000000000000000","111111111111101110","000000000000010101","111111111111101001","111111111111111110","111111111110101001","111111111110110001","000000000000000000","111111111111111001","000000000000100100","111111111111100010","000000000000001100","111111111111110100","000000000000000100","000000000000000011","111111111111110001","111111111111110010","111111111111111111","111111111111100101","111111111111100101","000000000000011000","111111111111110100","000000000000000001","000000000000010001","111111111111101111","111111111111111000","000000000000000000","000000000000001101","111111111111110000","111111111111110000","000000000000101011","000000000000000001","000000000000010101","111111111111110000","111111111111111110","111111111111111101","000000000000011101","000000000000000111","000000000000011011","000000000000011010","000000000000001111","000000000000010111","111111111111001001","000000000000001111","000000000000011001","000000000001000100","111111111111111010","111111111111110101","111111111111111000","111111111111111111","000000000000010011","000000000000000011","111111111111111010","000000000000001111","000000000000010010","111111111111101000","000000000000001101","111111111111110001","000000000000010011","111111111111110110","000000000000000010","111111111111101010","000000000000010000","111111111111110000","000000000000001010","111111111111101011","111111111111101010","000000000000101110","111111111111100110","000000000000001101","000000000000001000","000000000000010010"),
("111111111111111000","000000000000011111","000000000000010010","111111111111101011","111111111111101110","111111111111111100","111111111111110110","111111111111101100","000000000000000101","000000000000110001","000000000000000000","000000000000000111","111111111111110001","111111111111110010","000000000000000000","111111111111001101","111111111111011010","111111111111011111","000000000000000111","111111111111011100","000000000000010000","000000000000100000","111111111111111100","111111111111111100","111111111111111110","111111111111100010","000000000000011101","111111111111011100","111111111111111001","111111111111100000","111111111111111001","000000000000000001","111111111111110110","000000000000010110","000000000000000101","111111111111101111","000000000000001011","111111111111100000","000000000000001001","000000000000001010","000000000000010111","000000000000000001","111111111111110101","111111111111111111","000000000000000000","111111111111111011","000000000000001000","000000000000000110","000000000000100100","111111111111111001","111111111111100101","111111111111110001","000000000000001010","111111111111111110","111111111111101110","000000000000000111","000000000000000011","111111111111111010","000000000000100010","111111111111110111","000000000000000010","111111111110110101","111111111110111001","000000000000001010","000000000000011100","111111111111111110","111111111111010110","000000000000001000","111111111111000101","000000000000011110","111111111111110010","111111111111111000","111111111111111000","000000000000000011","000000000000001111","111111111111100000","111111111111110100","111111111111011110","000000000000100001","000000000000000111","000000000000001000","000000000000000011","000000000000001101","111111111111101011","111111111111111001","111111111111111111","000000000000011000","111111111111110110","000000000000011101","000000000000000110","000000000000010101","111111111111111000","000000000000001101","111111111111110101","000000000000010111","000000000000000111","000000000000011101","000000000000000100","111111111111010100","000000000000010011","111111111111110100","000000000000100111","000000000000001100","111111111111100111","111111111111101101","111111111111011111","000000000000010000","000000000000001001","111111111111100010","000000000000000000","000000000000011101","111111111111110100","111111111111101111","111111111111110110","000000000000000101","000000000000000111","111111111111111001","000000000000001011","000000000000000001","111111111111011100","000000000000000000","111111111111111110","000000000000000010","000000000001000100","000000000000000001","000000000000001000","111111111111101111","000000000000010011"),
("000000000000010110","111111111111100111","000000000000010001","000000000000000110","111111111111011010","111111111111110100","111111111111101011","000000000000100010","111111111111111101","000000000001010010","111111111111110111","000000000000100101","111111111111101000","111111111111111110","000000000000011111","111111111111010101","111111111111011011","111111111111110001","111111111111111111","111111111111011101","000000000000100110","000000000000000110","000000000000000100","111111111111111111","000000000000100011","111111111111101010","000000000000100000","111111111111110001","111111111111100010","111111111111111111","111111111111111010","111111111111100001","000000000000010000","000000000000000000","000000000000000111","111111111111110010","000000000000000101","111111111111101001","000000000000001001","000000000000010100","000000000000010110","000000000000001101","000000000000001000","000000000000000100","000000000000100001","000000000000000000","111111111111110100","000000000000001100","000000000000011101","111111111111110110","111111111111111010","000000000000000000","000000000000010101","111111111111110110","000000000000010110","000000000000011011","000000000000001011","111111111111110011","000000000000000101","000000000000001000","000000000000001111","111111111110111101","111111111111101100","000000000000000011","000000000000000110","000000000000001010","111111111111100011","111111111111101100","111111111111001000","000000000000000111","111111111111101100","111111111111011010","000000000000001000","111111111111110111","111111111111110010","111111111111111101","111111111111110101","111111111111110111","000000000000010111","000000000000001011","000000000000001110","000000000000000110","111111111111111000","111111111111000101","111111111111101011","000000000000011100","000000000000101000","111111111111110101","000000000000001110","000000000000011010","000000000000001001","000000000000000001","000000000000010010","000000000000000001","000000000000000100","000000000000000010","000000000000101111","111111111111111110","111111111111100100","111111111111011111","111111111111110101","000000000000001100","111111111111110110","000000000000000111","000000000000000100","111111111111100110","111111111111111110","111111111111110111","111111111111100010","000000000000000001","000000000000000101","111111111111011011","000000000000010000","000000000000001111","111111111111111111","000000000000000001","111111111111110100","000000000000001000","111111111111110010","111111111111111000","111111111111100010","000000000000000100","000000000000001001","000000000001010101","111111111111111101","000000000000000111","111111111111011110","000000000000000001"),
("000000000000000000","111111111111011111","000000000000000000","111111111111011110","111111111111001000","111111111111110000","000000000000000110","000000000000001010","111111111111110110","000000000001000111","111111111111100101","000000000000000000","111111111111010100","111111111111111010","111111111111100111","111111111111010101","111111111111101111","111111111111000100","111111111111011010","111111111111111000","000000000000000110","000000000000000001","111111111111110111","000000000000100000","111111111111111111","000000000000010100","000000000000101011","111111111111101101","111111111111100101","000000000000000111","000000000000001011","111111111111101010","111111111111111001","000000000000010001","000000000000001100","000000000000010111","000000000000000011","111111111111111001","111111111111111000","111111111111111101","111111111111111001","000000000000010101","111111111111111010","000000000000000101","000000000000100011","000000000000101111","111111111111101101","111111111111111111","000000000000000000","000000000000001110","000000000000010010","000000000000011000","111111111111101001","111111111111111011","111111111111111111","000000000000011111","000000000000011001","111111111111111111","000000000000010011","000000000000001000","000000000000010111","111111111111000101","111111111111101110","111111111111110001","000000000000001110","000000000000011001","000000000000001100","111111111111110101","111111111110011101","000000000000101101","000000000000000000","111111111111110101","111111111111110110","000000000000000001","000000000000011011","000000000000100010","000000000000001111","111111111111010000","000000000000001000","000000000000001111","000000000000000010","000000000000001010","000000000000001011","111111111110001100","111111111111101111","000000000000110010","000000000000001010","111111111111111101","000000000000010100","000000000000001101","000000000000001011","000000000000010111","000000000000010000","000000000000001001","000000000000010111","111111111111110001","000000000000011111","111111111111111010","000000000000011101","111111111111110100","111111111111100100","000000000000001000","111111111111111100","000000000000000111","000000000000100010","111111111111110011","000000000000000110","000000000000000000","111111111111011110","000000000000100100","000000000000001011","111111111111011001","000000000000011001","000000000000100101","111111111111011000","111111111111101101","111111111111110111","000000000000001001","000000000000010111","111111111111110001","111111111111011010","000000000000100101","111111111111111010","000000000000111011","000000000000101000","111111111111110100","111111111111010101","000000000000000111"),
("111111111111101101","111111111111010000","000000000000001011","111111111111100000","111111111111110100","111111111111101110","111111111111101001","000000000000000101","111111111111110111","000000000000101010","111111111111001011","111111111111110000","000000000000000100","111111111111111011","111111111111001110","111111111111001111","111111111111101001","111111111111100011","111111111111110011","111111111111110101","000000000000111010","111111111111110101","111111111111001010","000000000000010011","000000000000010100","000000000000000101","111111111111101101","111111111111001000","111111111111111110","000000000000100011","111111111111110111","000000000000000100","111111111111110101","000000000000001010","000000000000000100","000000000000000101","111111111111111011","000000000000010110","111111111111100010","000000000000001000","000000000000001011","000000000000100000","000000000000010011","000000000000010100","111111111111111111","000000000000100100","000000000000010011","111111111111011010","000000000000101001","000000000000100001","000000000000001100","111111111111100110","000000000000000101","000000000000111011","111111111111100111","111111111111111111","000000000000010000","000000000000010100","000000000000010100","000000000000000110","000000000000110000","111111111110110100","111111111111101110","111111111111110001","000000000000100010","111111111111111011","000000000000001001","000000000000001111","111111111110110000","111111111111110110","000000000000010110","111111111111101000","000000000000101000","000000000000001100","000000000000010110","000000000000101110","111111111111110011","111111111111001011","000000000000001000","111111111111110101","000000000000001100","111111111111100101","111111111111010111","111111111110100001","000000000000001010","000000000000011101","111111111111111110","000000000000001101","111111111111110100","000000000000110000","111111111111111011","000000000000100101","000000000000000000","000000000000010111","111111111111111100","111111111111111010","000000000000100101","111111111111110110","000000000000100011","111111111111110000","111111111111100010","111111111111100110","000000000000000111","000000000000011100","000000000000101101","000000000000001010","000000000000010101","111111111111100110","111111111111011110","000000000000001010","000000000000011001","111111111111001101","000000000000010011","000000000000100000","111111111111001010","000000000000000000","000000000000001100","000000000000001011","000000000000001010","111111111111110111","111111111111001111","000000000000011000","000000000000000001","000000000000001100","000000000000101011","000000000000000101","111111111111011100","000000000000010111"),
("111111111111101100","111111111111011110","111111111111110000","000000000000001010","000000000000001101","000000000000000000","111111111111100001","111111111111110001","000000000000000000","111111111111010110","111111111111011011","111111111111110111","000000000000000100","000000000000101110","111111111111010110","111111111111010111","111111111111110011","111111111111101110","111111111111110011","111111111111111100","000000000001010000","000000000000010101","111111111111000110","000000000000110100","111111111111101101","000000000000011111","111111111111010000","111111111111001110","000000000000011011","000000000000010101","000000000000000000","000000000000001111","111111111111110101","111111111111110101","000000000000011100","000000000000100101","111111111111110001","000000000000010100","111111111111100000","111111111111111000","111111111111100000","000000000000100001","000000000000100000","000000000000001101","111111111111111110","000000000000010111","000000000000011000","111111111111100000","000000000000011001","000000000000101001","000000000000011010","111111111111110000","000000000000010010","000000000000110000","000000000000000010","111111111111111100","000000000000100001","000000000000010110","111111111111111101","000000000000000111","000000000000011110","111111111111010101","111111111111100101","111111111111100010","000000000001001000","000000000000000001","000000000000100111","000000000000000001","111111111111011111","111111111111000111","000000000000000011","111111111111110111","000000000000111000","000000000000100100","000000000000100000","000000000000011011","000000000000000101","111111111111001011","000000000000000001","111111111111101111","000000000000000011","111111111111011101","111111111111010000","000000000000000000","000000000000011000","000000000000010100","111111111111100011","111111111111111100","111111111111011010","000000000000011010","111111111111110010","111111111111111000","000000000000101001","000000000000011110","000000000000000000","000000000000000110","000000000000110010","111111111111110010","000000000000010101","111111111111011100","111111111111100111","111111111111001100","000000000000011111","000000000000011101","000000000000011100","111111111111110110","000000000000100111","111111111111011111","111111111111100011","111111111111101001","000000000000100100","111111111111001100","000000000000001000","000000000000010111","111111111111010001","111111111111101111","000000000000010000","111111111111110101","111111111111111001","111111111111110000","111111111111000111","111111111111101010","000000000000011001","111111111111000111","000000000000010101","111111111111110011","111111111111100101","000000000000000101"),
("111111111111010010","111111111111011101","000000000000000100","111111111111110010","000000000000110110","111111111111111000","111111111111100010","111111111111011011","000000000000011110","111111111111001011","111111111111101010","111111111111101011","111111111111111000","000000000000011011","111111111111110111","111111111111011110","000000000000000100","000000000000000101","000000000000000001","111111111111010011","000000000000010011","000000000000001001","111111111111100001","000000000000000000","000000000000001100","000000000000000101","111111111111101101","111111111111110100","000000000000110000","111111111111110011","000000000000010111","000000000000001100","111111111111111010","111111111111100100","000000000000000111","000000000000100010","111111111111101011","000000000000011011","111111111111101100","000000000000000000","111111111111001011","000000000000101000","000000000000001101","000000000000011111","000000000000001100","000000000000011000","000000000000001111","111111111111101001","000000000000010001","000000000000001101","000000000000000011","111111111111100111","111111111111110000","111111111111111000","111111111111111111","000000000000011001","000000000000010100","000000000000000111","000000000000000001","000000000000000100","000000000000011000","000000000000001100","111111111111111011","000000000000001101","000000000000110000","111111111111111101","000000000000011110","111111111111101000","111111111111110100","111111111111011110","111111111111111110","000000000000000000","000000000000101101","000000000000101110","000000000000100100","000000000000000000","000000000000000000","111111111111100101","000000000000010010","111111111111111011","111111111111011111","111111111111111101","111111111111011011","000000000000110101","111111111111111101","000000000000000000","111111111111100001","000000000000000111","111111111111100010","000000000000011010","111111111111101001","111111111111111110","000000000000110011","111111111111111100","000000000000010001","000000000000000000","111111111111110100","111111111111100101","000000000000010111","111111111111011011","111111111111010010","111111111111100001","000000000000000010","111111111111110000","000000000000000000","111111111111100111","000000000000010010","111111111111100001","000000000000000011","111111111111111101","000000000000000001","111111111111100110","111111111111111111","000000000000010011","111111111111110011","111111111111011110","111111111111101001","111111111111111101","111111111111111111","111111111111110111","111111111111000000","111111111111111001","000000000000101101","111111111111011101","000000000000001101","111111111111010011","111111111111100011","000000000000001010"),
("111111111111001110","000000000000000010","000000000000011111","111111111111110111","000000000000010011","111111111111101101","111111111111100100","111111111111111001","000000000000010110","111111111111110110","111111111111101111","111111111111101011","000000000000001001","000000000000011011","000000000000001101","111111111111100110","000000000000100110","111111111111100011","000000000000001001","111111111111101110","000000000000001000","111111111111111100","000000000000010000","000000000000011101","000000000000001011","000000000000000110","111111111111101111","111111111111111011","000000000000010000","111111111111001101","111111111111110100","000000000000001111","111111111111110111","111111111111011010","000000000000000110","000000000000010001","111111111111111111","000000000000001010","111111111111111010","000000000000001001","111111111111011101","000000000000010001","000000000000011101","000000000000100000","000000000000000001","111111111111110110","111111111111110100","111111111111111000","000000000000001010","000000000000011000","000000000000001111","111111111111110010","111111111111101101","000000000000000100","000000000000011101","111111111111110111","111111111111111111","111111111111101011","000000000000001100","111111111111101111","000000000000001110","000000000000011011","111111111111111011","000000000000001011","000000000000011100","111111111111111010","000000000000001010","111111111111100100","111111111111110100","111111111111011111","111111111111111010","111111111111011001","000000000000000011","111111111111111100","000000000000010001","000000000000000101","000000000000010010","111111111111011111","000000000000010100","000000000000000100","111111111111100111","111111111111101110","111111111111101011","000000000000010011","000000000000000110","000000000000010000","111111111111110101","000000000000011010","111111111111100000","111111111111100110","111111111111101110","111111111111110011","000000000000111010","111111111111001101","000000000000100110","000000000000000011","111111111111110101","111111111111111100","000000000000000000","111111111111110110","111111111111110110","111111111111100000","111111111111101101","000000000000000111","111111111111111101","111111111111100000","000000000000001000","111111111111100011","000000000000010101","111111111111101011","000000000000010010","111111111111110000","111111111111110111","000000000000010001","111111111111101000","111111111111010111","000000000000000010","111111111111100000","111111111111111000","111111111111110011","111111111111101100","111111111111100010","000000000000010001","111111111111101000","000000000000011010","111111111111101000","111111111111010111","000000000000011001"),
("111111111110110010","000000000000000000","000000000000000011","111111111111111000","000000000000001110","111111111111101111","000000000000000010","000000000000000011","000000000000001100","000000000000000101","111111111111110000","111111111111101001","000000000000010101","000000000000100001","000000000000000110","111111111111110111","000000000000011111","111111111111110111","111111111111110110","000000000000001111","111111111111110111","000000000000010001","000000000000100100","111111111111110111","000000000000001001","000000000000000011","111111111111110111","000000000000000110","000000000000001010","111111111111010101","000000000000001011","000000000000011100","000000000000000001","111111111111110110","111111111111100111","000000000000011101","111111111111101101","111111111111111000","111111111111111011","111111111111111001","111111111111110101","000000000000000000","000000000000010101","000000000000001100","111111111111111000","000000000000000111","111111111111110101","111111111111111000","000000000000010101","000000000000101000","111111111111111011","111111111111110011","000000000000001100","111111111111111100","000000000000000100","000000000000001001","000000000000001101","000000000000001111","000000000000010000","111111111111110001","000000000000001110","000000000000100100","000000000000011000","000000000000010011","000000000000100011","111111111111111101","000000000000001000","000000000000001001","111111111111110111","000000000000000001","000000000000011000","000000000000000110","000000000000001111","000000000000101010","000000000000001100","000000000000000010","111111111111101010","000000000000000110","000000000000010001","000000000000001011","111111111111111101","000000000000010000","000000000000001010","000000000000010101","000000000000001100","000000000000010100","111111111111111000","000000000000001010","111111111111010000","111111111111011011","111111111111110110","000000000000010010","000000000000111111","111111111111001100","000000000000010001","000000000000000010","111111111111011011","000000000000001000","111111111111110011","000000000000101100","111111111111101010","111111111111100001","111111111111111001","000000000000001001","111111111111111010","000000000000000000","000000000000001101","000000000000000011","000000000000100100","111111111111110000","000000000000001010","000000000000001000","111111111111111011","111111111111111011","000000000000001101","111111111111001110","000000000000001000","111111111111111101","000000000000011101","000000000000010011","111111111111100111","111111111111100011","000000000000100110","000000000000011111","000000000000000111","111111111111111001","111111111111100110","000000000000001010"),
("111111111110111100","000000000000001101","111111111111111011","000000000000001111","111111111111011110","111111111111110000","000000000000000010","000000000000010011","000000000000000010","000000000000001011","000000000000000101","111111111111110110","000000000000000100","000000000000100111","111111111111111100","111111111111100101","000000000000000111","111111111111100111","000000000000000001","000000000000001011","000000000000001111","111111111111111101","000000000000011100","000000000000000000","111111111111110011","111111111111110010","000000000000001000","000000000000011010","111111111111101101","111111111111101101","111111111111101111","000000000000100010","000000000000010010","111111111111110001","111111111111101011","000000000000011101","111111111111111100","111111111111111100","000000000000000001","111111111111110010","000000000000001111","000000000000000010","000000000000010010","000000000000010010","000000000000000011","111111111111110001","111111111111111010","111111111111111100","111111111111111000","000000000000010100","111111111111100000","000000000000000100","111111111111111001","000000000000001111","000000000000010011","000000000000001000","111111111111100101","111111111111111000","000000000000001010","111111111111111010","111111111111110100","000000000000001111","000000000000000111","000000000000011111","000000000000011010","000000000000001010","000000000000011001","111111111111111100","111111111111101000","000000000000101010","000000000000000010","000000000000010001","111111111111110100","000000000000010000","000000000000000101","000000000000000010","111111111111110110","000000000000010101","111111111111101111","111111111111101111","111111111111110011","000000000000011001","111111111111101011","111111111111111110","000000000000000010","000000000000010101","000000000000000001","000000000000000000","111111111111100111","111111111111100100","111111111111101100","000000000000000110","000000000001001110","111111111111100001","000000000000011010","000000000000010001","111111111111011010","000000000000010001","000000000000001101","000000000000100001","111111111111011110","111111111111111110","111111111111110011","111111111111111001","000000000000001110","000000000000001100","111111111111111101","000000000000010101","000000000000010101","000000000000000000","000000000000001101","000000000000001010","111111111111100100","111111111111111011","000000000000010111","111111111111110010","111111111111101110","000000000000001001","111111111111111110","111111111111110100","111111111111011100","111111111111100111","111111111111110011","000000000000010010","000000000000001000","000000000000001111","111111111111010000","000000000000010101"),
("111111111110101001","111111111111011110","111111111111100000","000000000000011100","111111111111001111","000000000000010110","000000000000011100","111111111111111001","000000000000001001","111111111111111101","000000000000001111","000000000000000000","000000000000000011","000000000000011001","000000000000010110","111111111111110100","111111111111111101","000000000000001001","000000000000000100","000000000000010011","000000000000000000","000000000000001100","000000000000011010","111111111111110111","111111111111101011","000000000000001111","000000000000100001","000000000000100111","111111111111100111","111111111111101011","111111111111110110","000000000000100100","000000000000000100","111111111111100010","111111111111101100","000000000000011011","111111111111101100","111111111111111111","111111111111110110","000000000000000100","111111111111110001","000000000000000000","111111111111101101","000000000000010110","111111111111111100","111111111111100001","111111111111101011","111111111111101111","111111111111110111","000000000000001001","111111111111110111","000000000000011100","111111111111111111","111111111111110000","111111111111110011","111111111111111101","111111111111010100","000000000000000011","000000000000010010","111111111111111101","111111111111101010","111111111111110111","000000000000010101","000000000000001001","111111111111100111","111111111111111100","000000000000000001","000000000000000110","111111111111100001","000000000000011110","000000000000000100","111111111111101111","111111111111111110","111111111111111100","111111111111101001","111111111111100111","111111111111110110","000000000000001110","111111111111111110","111111111111111110","000000000000000110","000000000000000000","000000000000010110","111111111111100111","000000000000011001","000000000000011101","000000000000001110","111111111111111011","000000000000001100","111111111111101111","111111111111100000","000000000000000011","000000000000100101","111111111111111101","000000000000000011","000000000000010011","111111111110110101","000000000000000011","000000000000010110","000000000000101011","000000000000010001","111111111111101010","111111111111110100","000000000000001001","111111111111111010","000000000000000011","000000000000010011","000000000000010101","000000000000011010","000000000000001011","000000000000011011","000000000000010010","000000000000001001","000000000000001011","000000000000100000","000000000000001101","000000000000000101","000000000000001110","000000000000010000","000000000000001011","111111111111001010","000000000000000010","111111111111100110","000000000000010000","000000000000011111","111111111111110010","111111111111100100","000000000000001001"),
("111111111110111100","000000000000000000","000000000000001000","000000000000011110","111111111111011101","111111111111101111","000000000000011011","111111111111110110","000000000000001001","000000000000001101","111111111111110101","111111111111100111","111111111111110000","000000000000100001","000000000000000011","000000000000000010","111111111111100010","000000000000001001","111111111111101011","000000000000000101","000000000000010001","000000000000100100","000000000000001110","111111111111111001","000000000000001000","000000000000001110","000000000000010001","000000000000100101","111111111111010110","111111111111011010","111111111111100110","000000000000101000","000000000000010101","111111111111100101","111111111111110101","000000000000000001","111111111111110101","111111111111101111","000000000000000010","111111111111101001","111111111111100110","000000000000011011","111111111111101111","000000000000010001","111111111111101111","111111111111110110","000000000000000101","111111111111100001","111111111111100110","000000000000010001","000000000000001110","111111111111101111","000000000000010011","111111111111111100","111111111111011000","000000000000011100","111111111111110001","000000000000011101","000000000000100111","000000000000010001","111111111111110111","000000000000000010","000000000000100101","111111111111111011","111111111111011100","000000000000000100","111111111111110100","111111111111101111","111111111111010111","111111111111111111","000000000000010011","000000000000010010","000000000000010100","000000000000000110","000000000000000010","111111111111110101","111111111111111000","000000000000010000","111111111111111110","111111111111111010","111111111111100011","000000000000011110","111111111111111000","111111111111101010","000000000000001101","000000000000001110","000000000000000000","111111111111100100","000000000000010000","000000000000000011","111111111111101100","000000000000001100","000000000000101111","000000000000000101","000000000000000001","000000000000011000","111111111111100011","000000000000000111","111111111111110100","000000000000101111","000000000000000100","111111111111101100","000000000000000011","000000000000010101","111111111111110001","000000000000000111","000000000000001001","000000000000101001","000000000000010111","000000000000001100","000000000000000000","000000000000100010","111111111111100101","111111111111111111","000000000000011111","000000000000011101","000000000000010001","111111111111111001","000000000000010001","000000000000001111","111111111110110010","111111111111110001","111111111111110010","000000000000001100","000000000000010110","111111111111101101","111111111111011011","000000000000000110"),
("111111111110110111","000000000000000011","111111111111101100","000000000000010101","111111111111100011","111111111111110111","000000000000100000","111111111111010100","111111111111111010","111111111111110010","111111111111111111","111111111111111101","111111111111100110","000000000000000011","000000000000011000","111111111111110010","111111111111010110","111111111111110010","000000000000000001","111111111111110001","000000000000011101","000000000000110011","111111111111111011","111111111111111011","000000000000010000","000000000000000101","111111111111110000","000000000000000000","111111111111011101","111111111111101110","111111111111101011","000000000000011010","000000000000001000","111111111111000101","000000000000000001","111111111111101001","111111111111010110","111111111111010000","111111111111111000","111111111111010000","111111111111101101","111111111111101100","111111111111111000","111111111111100111","000000000000000011","111111111111010101","000000000000011010","111111111111111011","111111111111110010","000000000000010100","000000000000010001","111111111111111000","000000000000011011","000000000000000101","111111111111000011","000000000000010001","111111111111101111","000000000000010000","000000000000010011","111111111111101110","000000000000010010","111111111111110001","000000000000000000","111111111111111111","111111111111110110","000000000000000010","000000000000001110","111111111111111101","111111111111101001","000000000000000000","000000000000001101","000000000000000011","000000000000001011","111111111111110000","111111111111111110","111111111111100100","000000000000000111","000000000000101110","000000000000000010","000000000000010000","000000000000000010","000000000000001001","000000000000000111","000000000000001000","111111111111111010","111111111111111011","111111111111110111","111111111111011010","111111111111111111","111111111111111101","111111111111101101","000000000000000000","000000000000101010","000000000000010010","111111111111110101","111111111111111000","111111111111110110","000000000000000000","111111111111011011","000000000000011111","000000000000000101","111111111111111111","000000000000001101","111111111111110110","111111111111111001","111111111111111111","000000000000001011","000000000000010101","000000000000011110","000000000000001010","111111111111111011","000000000000100000","111111111111110001","000000000000001101","000000000000010011","000000000000010011","111111111111101110","111111111111110100","000000000000001000","111111111111100011","111111111110110101","000000000000000000","000000000000000100","000000000000001001","000000000000001111","111111111111011100","111111111111100001","000000000000001000"),
("111111111110010101","111111111111101011","111111111111111010","000000000000000100","111111111111100001","111111111111110110","000000000000000110","111111111111110001","111111111111111100","000000000000000000","111111111111101100","111111111111100100","000000000000010000","111111111111100000","000000000000010011","111111111111110110","111111111111110100","111111111111111101","000000000000010100","111111111111111010","000000000000110100","000000000000110101","000000000000010101","000000000000100101","000000000000000010","000000000000001001","000000000000000000","000000000000000000","111111111111101100","111111111111111010","111111111111011010","000000000000100000","000000000000001001","111111111110110010","000000000000000101","111111111111101111","111111111111011000","111111111110111001","000000000000010101","111111111111100001","111111111111101000","000000000000000111","111111111111111111","111111111111000101","111111111111111100","111111111111011001","111111111111110001","111111111111101001","111111111111111110","000000000000000000","000000000000001111","111111111111110111","000000000000000011","000000000000011001","111111111111100001","111111111111111100","111111111111010110","000000000000110000","000000000000100010","111111111111111100","000000000000000001","111111111111111011","111111111111101011","111111111111101110","111111111111011001","111111111111101110","000000000000011111","000000000000000000","111111111111110000","000000000000000101","000000000000001111","111111111111111000","000000000000011111","111111111111001111","111111111111110100","111111111111100101","000000000000000000","000000000000001001","000000000000100011","000000000000000111","111111111111101010","111111111111110101","000000000000000100","000000000000001000","111111111111111110","111111111111100111","000000000000000110","111111111111001111","111111111111011111","000000000000000010","111111111111110000","111111111111101110","000000000001000101","111111111111111111","000000000000010010","111111111111111000","111111111111110000","000000000000011011","111111111111110010","000000000000011010","111111111111110010","000000000000001100","000000000000001111","111111111111111111","000000000000000000","000000000000010101","111111111111111110","000000000000010001","000000000000010101","111111111111101100","000000000000001001","000000000000011100","111111111111011001","000000000000001010","000000000000010111","000000000000010000","000000000000000000","111111111111110000","000000000000010111","000000000000000000","111111111110110000","000000000000001000","111111111111100110","000000000000000000","000000000000001011","111111111111110001","111111111111100111","111111111111110111"),
("111111111110100011","000000000000000011","111111111111110111","111111111111111010","000000000000000000","111111111111110111","111111111111111100","111111111111111101","000000000000000110","000000000000011110","111111111111101110","111111111111111110","000000000000010100","111111111111110101","000000000000001000","111111111111110010","111111111111001001","000000000000011001","000000000000010100","111111111111011011","000000000000100111","000000000000010100","111111111111111110","000000000000100111","000000000000010110","111111111111111110","000000000000001100","000000000000000000","111111111111101011","000000000000000111","111111111111100010","000000000000100100","000000000000011011","111111111111011111","000000000000000000","111111111111011010","111111111111101001","111111111111100100","000000000000000110","111111111111100000","111111111111110100","000000000000001010","111111111111010000","111111111111000111","111111111111110100","111111111111100011","000000000000001110","111111111111110111","111111111111111100","000000000000000010","111111111111111011","000000000000000000","000000000000011101","000000000000001010","111111111111011100","000000000000000000","000000000000000000","000000000000000000","000000000000011000","111111111111111011","000000000000001011","111111111111100001","111111111111001101","111111111111101001","111111111111011111","111111111111110101","000000000000101010","000000000000100000","111111111111110010","000000000000001000","111111111111111010","111111111111100010","000000000000011010","111111111111100000","000000000000000011","111111111111101101","111111111111101101","000000000000010110","111111111111110010","000000000000001010","111111111111110110","000000000000010111","111111111111011100","111111111111011000","111111111111111011","111111111111010101","111111111111110000","111111111111001010","111111111111110111","111111111111111000","111111111111011111","000000000000000000","000000000000110110","000000000000011100","111111111111111011","000000000000011010","111111111111111101","000000000000010001","111111111111111111","111111111111010000","000000000000000100","000000000000010100","000000000000000111","111111111111111100","000000000000110011","000000000000010011","111111111111111101","000000000000000000","111111111111101100","111111111111011100","000000000000000000","000000000000001011","111111111111111110","111111111111110001","111111111111111010","000000000000001110","000000000000000111","111111111111110010","000000000001001000","111111111111111011","111111111110011111","000000000000010110","111111111111110101","111111111111110010","111111111111110000","111111111111100000","111111111111011101","000000000000001100"),
("111111111111001101","000000000000010010","111111111111101001","111111111111011111","111111111111000101","111111111111111001","111111111111110011","111111111111111101","111111111111111101","000000000000001010","000000000000000000","000000000000101100","000000000000001110","000000000000001111","111111111111100111","000000000000011011","111111111110111001","000000000000011101","000000000000010100","111111111111111101","000000000000101000","111111111111110001","000000000000001000","000000000000000001","000000000000111001","111111111111111011","000000000000000110","111111111111111111","111111111111111101","000000000000000011","000000000000010110","000000000000010000","000000000000010100","111111111111101010","000000000000011010","111111111111011101","111111111111100101","111111111111101111","000000000000110100","111111111111010010","000000000000000010","000000000000010100","111111111111000111","111111111111001001","111111111111111110","111111111111001010","000000000000000100","111111111111111111","000000000000001000","111111111111001100","000000000000011100","000000000000000110","000000000000111001","111111111111111101","111111111111001010","111111111111100011","000000000000011101","111111111111111011","111111111111111110","111111111111111000","000000000000001001","111111111111110110","111111111111000010","111111111111011000","111111111111010010","000000000000101000","000000000000011111","000000000000011111","111111111111011110","000000000000011110","000000000000010110","111111111111101110","000000000000110001","111111111111001000","000000000000000000","111111111111101100","000000000000011011","111111111111110001","111111111111011100","111111111111110110","000000000000001000","000000000000010011","111111111111000101","111111111111000000","000000000000000111","111111111111010001","111111111111110001","111111111111010011","111111111111100100","111111111110111000","111111111111000111","111111111111111111","000000000001101011","000000000000010010","111111111111101011","000000000000001101","000000000000010111","000000000000001100","111111111111111011","111111111111001111","000000000000100010","000000000000101010","000000000000001101","000000000000010101","000000000001000011","000000000000100010","111111111111101100","000000000000000011","111111111111011000","111111111111011100","000000000000001110","000000000000010100","000000000000010110","111111111111101000","000000000000000000","000000000000000000","000000000000011010","111111111111110010","000000000001001101","111111111111011110","111111111111001111","000000000000011100","111111111111011000","111111111111101010","111111111110111101","111111111111110010","000000000000000110","000000000000010100"),
("000000000000000110","111111111111110000","000000000000000000","000000000000010100","111111111111010110","000000000000000010","111111111111111100","000000000000011001","000000000000011001","111111111111110110","000000000000001001","000000000000001000","111111111111110001","000000000000010001","111111111111101001","000000000000000101","111111111110111111","000000000000100111","000000000000001010","000000000000000011","000000000001000010","111111111111101001","111111111111100010","111111111111111111","000000000000100010","000000000000011101","000000000000100111","111111111111101100","111111111111100010","111111111111101011","000000000000100111","111111111111101111","000000000000101011","111111111111110101","000000000000101011","111111111111101001","111111111111111000","111111111111111101","000000000000100010","111111111111110110","111111111111110001","000000000000001111","111111111111010110","111111111111011111","000000000000011101","111111111111010111","111111111111100000","000000000000000100","111111111111111001","111111111111001100","000000000000000010","000000000000001001","000000000000001011","000000000000000011","000000000000000111","000000000000010011","000000000000010111","111111111111110101","111111111110111101","111111111111110011","000000000000001010","111111111111100110","111111111111111101","111111111111001000","111111111111001011","111111111111110111","000000000000100100","111111111111111010","000000000000100010","000000000000001100","000000000000001011","000000000000001100","000000000000101010","111111111111101011","111111111111101011","000000000000100000","000000000000110100","111111111111101010","111111111111010010","111111111111100110","111111111111101100","000000000000110000","111111111111110010","111111111111011000","000000000000010001","111111111111001001","111111111111011110","111111111111110111","111111111111011101","111111111111110000","111111111111001011","000000000000001000","000000000000011010","111111111111000110","111111111111111010","111111111111101100","000000000000100110","000000000000100110","111111111111101111","111111111111110011","000000000000111000","111111111111111111","111111111111100000","000000000000010110","000000000000111000","000000000000000100","000000000000000000","111111111111100101","111111111111111101","111111111111010111","000000000000010000","000000000000001011","000000000000000010","111111111111111111","111111111111101001","111111111111110011","000000000000000100","000000000000011001","000000000000011111","111111111111110110","111111111111101010","000000000000011001","000000000000000010","111111111111000010","111111111111100110","111111111111011101","111111111111111111","000000000000010000"),
("111111111111110000","111111111111010001","000000000000001110","000000000000000001","111111111111011010","111111111111110001","111111111111111010","111111111111100010","000000000000010001","111111111111011110","000000000000001110","000000000000110001","111111111111110001","111111111111100101","111111111111001001","111111111111101000","111111111111100111","000000000000000011","111111111111111110","000000000000001010","000000000000100111","111111111111010000","111111111111100111","000000000000011001","000000000000011100","000000000000011010","000000000000101011","111111111111100010","111111111111110111","000000000000010010","000000000000111000","111111111111110101","000000000000100111","111111111111110111","000000000000111111","000000000000001001","111111111111111011","000000000000011000","000000000000001101","000000000000011000","000000000000010000","000000000000100101","111111111111011001","111111111111101010","000000000000110101","111111111111101011","111111111111101100","000000000000010101","000000000000100001","111111111111111111","000000000000101000","000000000001000000","000000000000010000","000000000000101111","111111111111101100","000000000000011100","000000000000010110","111111111111011010","111111111111101010","000000000000001100","000000000000111101","111111111111001111","111111111111110101","111111111111101101","111111111111100001","000000000000011101","000000000000011010","000000000000001000","111111111111111010","000000000000011100","000000000000001101","000000000000010100","000000000000000011","111111111111100011","000000000000000110","111111111111110101","000000000000011111","111111111111111001","111111111111110000","000000000000000010","000000000000010011","000000000000101000","111111111111100101","111111111111001011","000000000000000001","111111111110110110","000000000000000000","111111111111111111","111111111111111000","000000000000000010","111111111111100111","000000000000000001","000000000000100110","111111111111011111","000000000000000001","111111111111011111","000000000000000000","000000000000100000","111111111111110001","111111111111110110","111111111111110100","000000000000001100","111111111111101100","000000000000000101","000000000000110111","000000000000010111","000000000000001011","111111111111010110","111111111111110001","111111111110111101","000000000000010101","000000000000001100","000000000000001110","000000000000010110","000000000000010000","111111111111000110","111111111111110110","000000000000110001","000000000000101110","000000000000001011","111111111111110001","111111111111111010","111111111111011101","111111111111110000","111111111111001011","000000000000000100","000000000000010111","000000000000100101"),
("111111111111100101","000000000000100011","000000000000011000","111111111111111001","000000000000000111","111111111111101010","000000000000001110","111111111111100111","000000000000100001","000000000000001011","000000000000010001","000000000000010001","000000000000010001","111111111111110011","111111111111110000","111111111111110010","111111111111111011","000000000000000000","000000000000001101","111111111111100110","000000000000011011","000000000000010100","111111111111101011","111111111111111000","000000000000001110","000000000000000000","111111111111100100","111111111111100110","111111111111111011","000000000000010001","111111111111111110","000000000000000000","111111111111111000","111111111111101101","000000000000010111","111111111111101100","000000000000000010","111111111111111000","111111111111011111","000000000000011100","000000000000010000","000000000000101000","111111111111111010","111111111111111101","111111111111101011","000000000000000010","000000000000010001","111111111111110101","000000000000001001","111111111111101111","000000000000001011","000000000000000011","000000000000100001","000000000000010101","000000000000010001","000000000000011011","000000000000001111","111111111111111110","000000000000001111","000000000000001001","000000000000010010","000000000000001000","111111111111111111","111111111111100110","000000000000000100","111111111111111000","000000000000000000","111111111111110010","111111111111110001","000000000000001000","111111111111111010","000000000000000011","000000000000011000","111111111111110001","000000000000001110","000000000000001101","111111111111101010","000000000000001000","111111111111101100","111111111111111110","111111111111011100","111111111111111010","111111111111011011","000000000000001101","000000000000001000","111111111111101101","111111111111110101","111111111111110000","111111111111010100","000000000000010101","111111111111101110","000000000000001001","000000000000010011","111111111111101001","000000000000011001","111111111111111111","000000000000001011","000000000000000110","111111111111110101","000000000000011100","111111111111100100","111111111111101111","111111111111111100","000000000000000000","000000000000010101","111111111111111010","000000000000010110","000000000000000010","111111111111111110","000000000000001011","000000000000001001","000000000000000011","111111111111110101","111111111111100011","000000000000001101","111111111111100001","111111111111111001","000000000000001000","111111111111110101","000000000000000110","000000000000001000","111111111111101110","000000000000000000","000000000000000110","111111111111101100","111111111111110010","111111111111101011","000000000000001001"),
("111111111111110000","000000000000001001","000000000000010000","111111111111101111","000000000000011100","111111111111101100","000000000000000101","000000000000000001","111111111111101110","111111111111111010","111111111111101111","000000000000010011","111111111111110000","111111111111110010","000000000000000010","000000000000000100","000000000000000001","111111111111111011","000000000000100001","111111111111110011","000000000000100001","000000000000001110","000000000000000111","111111111111111001","000000000000001100","111111111111110011","000000000000010000","111111111111100111","000000000000011111","000000000000010011","000000000000000000","000000000000000010","111111111111110111","000000000000000111","111111111111110001","111111111111101010","000000000000100010","111111111111111011","000000000000010100","000000000000010001","000000000000100101","111111111111110110","111111111111111111","111111111111111111","111111111111101101","000000000000001110","111111111111110011","000000000000010010","000000000000100010","111111111111111111","111111111111101110","111111111111110000","000000000000001000","000000000000000111","000000000000010010","111111111111111110","111111111111111100","000000000000000011","000000000000011100","000000000000010010","111111111111111110","111111111111110010","111111111111110001","000000000000001101","000000000000001001","000000000000000101","000000000000001110","111111111111110101","000000000000001001","000000000000011000","111111111111011100","111111111111111001","111111111111111111","111111111111111101","111111111111101110","000000000000000111","111111111111101111","111111111111111000","000000000000000110","111111111111111111","000000000000001010","111111111111111001","000000000000000011","000000000000001011","000000000000000000","000000000000011010","000000000000011110","111111111111111001","111111111111110100","000000000000001111","000000000000000110","111111111111110010","111111111111110011","000000000000010000","000000000000010111","000000000000000101","111111111111111001","111111111111101000","000000000000001110","111111111111111111","000000000000001110","000000000000000100","111111111111111110","111111111111101001","000000000000000110","111111111111101001","111111111111111110","000000000000010010","000000000000100001","000000000000001000","111111111111111111","111111111111100010","111111111111110011","000000000000010111","000000000000001001","111111111111110000","111111111111011111","111111111111111011","000000000000001110","111111111111111011","000000000000010011","111111111111110110","111111111111110000","000000000000001111","000000000000010100","111111111111110101","000000000000010010","000000000000000010"),
("111111111111110010","000000000000001101","000000000000000011","111111111111110000","000000000000010000","000000000000000101","000000000000000101","111111111111101001","111111111111110001","111111111111111100","111111111111111111","000000000000000000","111111111111111100","000000000000010110","000000000000001101","111111111111101111","000000000000000000","000000000000000100","000000000000011011","000000000000011010","111111111111111100","000000000000111110","000000000000001100","000000000000000100","000000000000001100","111111111111101110","000000000000001111","111111111111110110","000000000000000001","000000000000011011","111111111111110110","000000000000001001","111111111111100110","000000000000001100","111111111111111111","111111111111101110","000000000000000111","000000000000001010","111111111111111010","000000000000000100","000000000000000000","000000000000001111","111111111111111001","111111111111111010","111111111111110100","000000000000001011","111111111111111100","111111111111110000","111111111111111111","000000000000000111","111111111111101110","000000000000000000","111111111111111010","000000000000001010","000000000000010011","000000000000000011","111111111111101100","000000000000001110","000000000000001011","000000000000001110","000000000000000111","000000000000000000","111111111111111000","111111111111111100","111111111111110000","000000000000000101","000000000000000100","111111111111101100","000000000000010101","111111111111111101","111111111111111110","000000000000000010","000000000000001100","000000000000000010","111111111111110101","000000000000000110","000000000000000100","000000000000000001","111111111111111101","111111111111111011","111111111111111101","111111111111110001","111111111111101000","111111111111111100","111111111111110100","111111111111111111","000000000000100001","111111111111110100","111111111111110001","000000000000001101","111111111111110111","111111111111100010","000000000000001001","000000000000000100","111111111111110101","111111111111111111","111111111111100010","111111111111100111","000000000000011000","000000000000011100","111111111111101011","111111111111111101","111111111111111110","000000000000000000","000000000000010011","111111111111110101","111111111111101110","000000000000001010","111111111111111001","111111111111110111","111111111111111101","111111111111001101","111111111111101010","000000000000001010","000000000000000001","000000000000000110","000000000000001000","111111111111111010","111111111111101010","111111111111111100","111111111111111001","111111111111110111","000000000000000100","000000000000100100","000000000000010101","111111111111101011","111111111111111100","111111111111110101"),
("111111111111111001","111111111111111111","000000000000000000","111111111111100100","000000000000010100","111111111111110100","111111111111110111","111111111111100000","111111111111111111","000000000000001010","000000000000011010","111111111111111110","000000000000011011","000000000000100110","000000000000001010","111111111111100100","111111111111110110","111111111111111010","000000000000011101","111111111111111010","000000000000100101","000000000000001000","000000000000000000","111111111111011100","000000000000010001","111111111111101000","000000000000001000","111111111111111011","000000000000101010","000000000000000111","111111111111101011","000000000000001100","111111111111100100","111111111111111100","000000000000010100","111111111111101101","000000000000001101","111111111111111110","111111111111110010","000000000000011110","000000000000101000","000000000000001100","000000000000011010","111111111111101000","111111111111101001","111111111111110011","111111111111110111","111111111111010110","000000000000100000","000000000000010110","111111111111011000","111111111111100111","000000000000001011","000000000000000000","000000000000000100","111111111111111100","111111111111100111","000000000000001001","000000000000001000","000000000000000000","111111111111111010","111111111111011010","111111111111100110","111111111111110001","000000000000010100","000000000000100001","000000000000011110","111111111111111100","111111111111100110","000000000000000110","111111111111011111","111111111111110111","000000000000010011","000000000000001001","111111111111101000","111111111111101101","111111111111100010","111111111111110110","000000000000000100","000000000000000100","111111111111110011","111111111111110100","000000000000000000","000000000000001111","111111111111011110","000000000000010000","000000000000011001","000000000000000100","111111111111110111","000000000000011011","000000000000010010","111111111111010010","000000000000010010","000000000000010110","000000000000010001","000000000000001001","111111111111110100","111111111111110111","111111111111111101","000000000000100101","111111111111110010","111111111111110011","000000000000000011","111111111111100001","000000000000010111","000000000000000110","111111111111100010","111111111111110100","111111111111011111","000000000000000000","000000000000010011","111111111111110101","111111111111011111","000000000000100011","111111111111111000","111111111111111101","111111111111100110","111111111111111001","111111111111101111","111111111111111110","000000000000010010","111111111111101111","000000000000001111","000000000000000011","000000000000010110","111111111111101010","000000000000000111","111111111111110111"),
("111111111111111010","000000000000001001","000000000000001010","111111111111111101","000000000000001110","111111111111111100","000000000000001011","000000000000011011","000000000000001011","000000000000100100","000000000000000001","000000000000001110","111111111111111100","000000000000011000","111111111111110000","111111111111100111","111111111111011001","111111111111110110","111111111111110101","111111111111100011","111111111111111101","000000000000000010","111111111111100100","111111111111101111","111111111111111010","111111111111110101","000000000000010100","111111111111111000","111111111111111011","111111111111101001","111111111111101110","000000000000000110","111111111111111101","111111111111101100","111111111111110111","111111111111101011","111111111111110111","000000000000010001","111111111111101010","000000000000000000","000000000000000111","000000000000000000","000000000000110000","000000000000001001","111111111111100001","111111111111110011","000000000000000011","111111111111111011","000000000000001011","000000000000110010","111111111111100111","111111111111110111","000000000000011111","000000000000001110","000000000000010010","000000000000001111","111111111111111001","111111111111111010","000000000000011101","111111111111101100","000000000000001001","111111111111000110","111111111111011111","111111111111011110","111111111111110011","000000000000000100","000000000000000111","111111111111101101","111111111111011000","000000000000010101","000000000000011001","000000000000000100","000000000000011101","000000000000010011","111111111111110010","111111111111101001","000000000000000010","111111111111100000","111111111111110111","111111111111110010","111111111111100011","000000000000001010","111111111111010001","111111111111111100","000000000000001000","111111111111110111","111111111111111111","111111111111100011","111111111111100001","000000000000000001","111111111111100000","111111111111111101","000000000000011001","111111111111110000","000000000000000110","111111111111111011","111111111111010010","111111111111110110","000000000000011010","000000000000010010","111111111111011010","111111111111110001","111111111111100011","111111111111111001","111111111111110110","000000000000010111","000000000000001111","000000000000010010","111111111111110001","111111111111100101","000000000000100000","000000000000010100","000000000000000001","000000000000011101","000000000000011010","111111111111011110","111111111111100011","000000000000000001","111111111111011010","000000000000010001","111111111111100010","111111111111101110","000000000000000101","000000000000001011","111111111111111010","000000000000001010","111111111111110000","000000000000000011"),
("000000000000011010","000000000000001101","111111111111101101","000000000000011000","111111111111100111","111111111111110010","111111111111111111","000000000000111010","111111111111101011","111111111111011111","000000000000110110","111111111111111100","111111111111010100","000000000000001000","111111111111110111","111111111111101000","111111111111100000","111111111111111111","111111111111110010","111111111111010101","000000000000001100","000000000000011000","111111111111111001","111111111111110100","000000000000010011","000000000000010000","111111111111110100","111111111111101110","111111111111111000","111111111111101110","000000000000001110","000000000000100010","000000000000000010","111111111111111000","111111111111110010","000000000000000101","111111111111110010","000000000000000100","111111111111010111","111111111111101111","000000000000011110","000000000000100000","000000000000011010","000000000000011101","000000000000001011","111111111111111011","000000000000000010","111111111111011011","000000000000000111","111111111111111111","111111111111000110","111111111111111110","000000000000010011","000000000000100010","111111111111110000","000000000000011110","111111111111011111","111111111111110110","000000000000010101","000000000000001100","000000000000110010","111111111110100011","111111111111010101","111111111111100001","111111111111100101","111111111111111011","000000000000000100","111111111111101110","111111111110111101","111111111111011111","000000000000010111","111111111111110011","000000000000010101","000000000000100001","000000000000001011","111111111111110110","111111111111110101","111111111111111010","111111111111100110","111111111111101001","111111111111110011","000000000000010001","111111111111011110","000000000000001001","000000000000001101","111111111111010101","000000000000101001","111111111111110110","111111111111000000","111111111111100100","111111111111010011","111111111111100101","000000000000001100","000000000000000010","000000000000011111","111111111111100010","111111111111000100","000000000000001101","000000000000011011","000000000000101001","111111111111111111","111111111111100111","000000000000001110","000000000000000010","000000000000001100","000000000000010101","000000000000001011","000000000000011010","111111111111101000","111111111111101100","000000000000001000","000000000000100000","111111111111110011","000000000000000011","000000000000000100","000000000000010100","111111111111111100","000000000000010011","111111111111011111","000000000000010001","111111111111101101","111111111111111000","000000000000001001","000000000000101011","111111111111011101","111111111111101010","111111111111010101","000000000000010101"),
("111111111111110110","000000000000000110","111111111111111110","000000000000001000","000000000000001011","111111111111111010","000000000000001101","000000000000001011","111111111111110111","000000000000000000","000000000000010101","000000000000000101","111111111111101011","111111111111011100","000000000000001101","111111111111011001","111111111111110001","111111111111111010","111111111111101001","111111111111100011","111111111111110111","000000000000101010","111111111111110100","111111111111101001","000000000000010000","000000000000010010","111111111111111101","111111111111100110","111111111111110111","000000000000000111","111111111111111101","000000000000000100","000000000000000101","111111111111011011","111111111111110010","111111111111110011","111111111111101000","111111111111111111","111111111111100110","111111111111110101","111111111111111010","000000000000000000","000000000000101000","111111111111110001","000000000000100000","111111111111100001","111111111111110011","111111111111100000","000000000000011010","000000000000001111","111111111111000110","111111111111110001","000000000000000000","000000000000001110","111111111111011001","000000000000010101","111111111111011111","111111111111011101","000000000000000011","000000000000001101","000000000000100000","111111111110101111","111111111111100000","000000000000000011","111111111111010001","000000000000001101","111111111111101010","111111111111111101","111111111111010011","000000000000000101","000000000000100010","111111111111101000","111111111111100100","000000000000001011","000000000000010101","111111111111110110","111111111111110101","111111111111100100","111111111111110101","111111111111100010","111111111111110010","000000000000010111","111111111111100010","111111111111010110","111111111111101010","111111111111010011","000000000000110000","111111111111110001","111111111111001110","111111111111111111","111111111111100111","111111111111101010","000000000000000111","111111111111011100","000000000000101101","111111111111101110","111111111111111111","000000000000001110","111111111111100011","000000000000000111","000000000000000011","000000000000001011","000000000000000110","111111111111111111","111111111111111111","000000000000000011","000000000000101100","000000000000000010","111111111111100110","111111111111101011","000000000000011010","000000000000000111","000000000000000101","000000000000000001","000000000000000011","111111111111111011","111111111111111111","000000000000010010","111111111111011110","111111111111101001","111111111111101011","111111111111101101","000000000000010001","000000000000110110","111111111111010010","111111111111110100","111111111111010110","000000000000001100"),
("000000000000000110","000000000000101110","000000000000001010","000000000000000100","000000000000001010","111111111111111011","000000000000011111","111111111111110001","111111111110111100","000000000000011111","000000000000011100","000000000000010001","111111111111101110","111111111111111110","111111111111110110","111111111111001111","111111111111101100","111111111111110010","111111111111101010","111111111111100001","000000000000001100","000000000000011000","000000000000100011","111111111111011110","000000000000010110","000000000000001001","000000000000000010","111111111111100011","111111111111100111","111111111111110111","000000000000001101","000000000000000000","111111111111111011","111111111111010011","111111111111100101","000000000000010001","111111111111111110","111111111111110000","000000000000010111","111111111111111000","000000000000011110","000000000000000111","111111111111110101","111111111111011111","000000000000011010","111111111111101110","111111111111111011","111111111111100101","000000000000010010","111111111111101110","111111111111111000","000000000000001000","000000000000000101","000000000000010010","111111111111010010","000000000000000110","111111111111110010","111111111111011001","000000000000011111","111111111111111110","111111111111111111","111111111110111101","111111111110111010","000000000000011100","111111111111010111","000000000000100011","111111111111100010","000000000000100100","111111111111100010","111111111111111101","000000000000000100","111111111111100001","111111111111100111","111111111111111011","000000000000001010","000000000000010001","111111111111101110","111111111111110010","111111111111111011","111111111111011100","000000000000000110","000000000000010111","111111111111101001","111111111111100010","000000000000000100","111111111111010100","000000000000101001","111111111111111000","111111111111110011","111111111111101011","111111111111101111","000000000000001010","111111111111111101","111111111111110101","000000000000000101","111111111111111011","000000000000001001","111111111111101001","111111111111010000","000000000000100000","000000000000010110","000000000000011100","111111111111101111","000000000000010000","111111111111101010","000000000000011101","000000000000010011","000000000000000110","000000000000000101","111111111111011111","000000000000000011","000000000000011010","000000000000000101","000000000000000101","000000000000001000","000000000000000000","000000000000010011","000000000000001010","000000000000000100","111111111111101100","111111111111101111","111111111111111011","000000000000001011","000000000000000011","111111111111011111","000000000000100110","111111111111100101","000000000000001111"),
("000000000000000011","000000000000001101","000000000000100101","000000000000000101","000000000000010010","000000000000001001","111111111111111100","111111111111101100","111111111111001001","000000000000010000","000000000000011010","000000000000010111","111111111111111101","111111111111110101","000000000000011110","111111111111010011","111111111111101011","111111111111111110","000000000000001010","111111111111001100","000000000000010001","000000000000001111","000000000000001010","111111111111100111","000000000000000001","111111111111111010","000000000000001000","111111111111110111","111111111111110100","111111111111100011","111111111111111101","000000000000000111","111111111111111100","111111111111100011","000000000000000010","111111111111110100","000000000000001000","111111111111110101","111111111111111011","000000000000000100","000000000000000010","000000000000001011","111111111111110111","111111111111100111","000000000000000110","000000000000000011","111111111111101101","111111111111101010","000000000000001100","111111111111101010","111111111111100111","111111111111111010","000000000000011010","000000000000000111","111111111111101010","000000000000000000","000000000000000000","111111111111100001","000000000000001000","000000000000001011","000000000000000101","111111111110011111","111111111111000011","000000000000000001","111111111111111100","000000000000001110","111111111111110001","000000000000011100","111111111110110101","000000000000000010","000000000000001010","111111111111011110","000000000000010100","000000000000010111","111111111111101001","000000000000010000","000000000000001011","111111111111101100","000000000000001011","111111111111100101","111111111111111011","111111111111111100","000000000000001011","111111111111101010","000000000000001010","000000000000000000","000000000000010011","111111111111110111","000000000000011000","111111111111110011","111111111111110011","000000000000001010","000000000000011100","111111111111111011","000000000000010011","111111111111101001","000000000000000000","000000000000001101","111111111111100100","000000000000010001","000000000000000110","000000000000001110","000000000000001100","000000000000011010","111111111111101100","000000000000010111","000000000000001010","000000000000001011","000000000000001110","111111111111111110","000000000000000010","000000000000000000","111111111111111101","111111111111101010","000000000000000111","111111111111101110","000000000000000001","000000000000011101","000000000000000011","111111111111100010","000000000000000011","111111111111111000","111111111111110111","000000000000100101","111111111111100100","000000000000001000","000000000000001000","111111111111110110"),
("111111111111111010","000000000000011100","000000000000011001","000000000000001101","000000000000100010","111111111111111001","111111111111110010","111111111111100010","111111111111011110","000000000000110110","000000000000011111","000000000000000110","111111111111011111","111111111111111101","000000000000101011","111111111111010010","111111111111010111","111111111111101011","000000000000010000","111111111111101010","000000000000000110","000000000000111000","111111111111111110","111111111111001101","000000000000001100","111111111111111101","111111111111111001","111111111111110111","111111111111110101","111111111111110001","111111111111101111","111111111111110011","000000000000000101","111111111111111100","000000000000000000","111111111111111011","111111111111110101","111111111111100001","000000000000001001","111111111111110100","111111111111111110","000000000000000011","111111111111111100","111111111111110000","000000000000000010","000000000000000010","000000000000001010","111111111111111001","000000000000010110","000000000000001000","111111111111011110","000000000000000110","111111111111111110","000000000000010101","111111111111110100","000000000000001110","111111111111110001","111111111111111100","000000000000001101","111111111111111111","111111111111110111","111111111110110100","111111111111010010","000000000000000110","111111111111110110","000000000000101100","111111111111010111","000000000000010100","111111111110101001","000000000000010101","111111111111100011","111111111111101100","000000000000010011","000000000000000000","111111111111101011","000000000000010101","000000000000000001","111111111111100111","000000000000000110","000000000000000000","111111111111110001","111111111111110010","000000000000000101","111111111111111011","111111111111100110","111111111111111001","000000000000100000","000000000000000000","000000000000011101","111111111111110001","111111111111110100","000000000000000001","000000000000001110","000000000000000110","000000000000010011","000000000000001100","000000000000010100","000000000000000101","111111111111100110","000000000000001001","000000000000100000","000000000000001100","111111111111110011","111111111111111100","111111111111110110","111111111111111000","000000000000000110","111111111111111100","111111111111111100","000000000000000001","000000000000001110","000000000000010011","111111111111110110","111111111111110011","111111111111111111","111111111111111101","111111111111111010","000000000000010011","000000000000010010","111111111111011101","111111111111110110","111111111111111111","111111111111111110","000000000000101011","111111111111101001","000000000000001111","000000000000000000","111111111111110101"),
("000000000000000111","000000000000001010","000000000000100111","000000000000001101","000000000000001111","000000000000011010","000000000000011000","111111111111110011","111111111111100001","000000000001011010","000000000000010000","000000000000010100","111111111111110010","000000000000000010","000000000000000000","111111111111011000","111111111111011101","000000000000000000","000000000000001100","111111111111100101","111111111111111010","000000000000100110","000000000000000110","111111111111110111","111111111111111010","111111111111111010","000000000000001100","111111111111111001","111111111111111101","000000000000010100","000000000000000110","111111111111101111","000000000000001011","000000000000011011","000000000000000010","111111111111111001","111111111111101111","111111111111111000","111111111111111001","000000000000001111","000000000000001100","000000000000000000","111111111111110100","000000000000000110","111111111111111101","000000000000000110","111111111111101101","000000000000000001","000000000000011001","111111111111110111","111111111111101010","000000000000001011","000000000000010100","111111111111111111","000000000000000010","000000000000001000","111111111111110000","111111111111110100","000000000000001111","111111111111110010","111111111111110111","111111111111001000","111111111110111110","000000000000011010","000000000000011100","000000000000000001","111111111111100101","000000000000011001","111111111110011010","000000000000001010","111111111111101001","111111111111011001","000000000000000100","000000000000000101","111111111111110010","000000000000000111","000000000000001111","111111111111110001","111111111111111010","000000000000001001","111111111111111011","000000000000001111","000000000000010110","111111111111000100","111111111111110110","111111111111111110","000000000000010100","000000000000010110","000000000000001110","000000000000001101","111111111111110101","111111111111111011","000000000000011000","000000000000010110","111111111111111111","000000000000010110","000000000000100001","000000000000001111","111111111111100010","111111111111111000","000000000000011111","000000000000101010","111111111111111110","000000000000000101","000000000000000001","111111111111110110","000000000000000010","111111111111111101","111111111111101001","000000000000010001","000000000000001010","111111111111110111","000000000000010011","111111111111110100","111111111111101000","000000000000000011","000000000000000000","000000000000001100","000000000000001101","111111111111100101","111111111111111111","111111111111011100","000000000000000100","000000000000101000","111111111111110111","000000000000000101","111111111111111010","000000000000000010"),
("000000000000010111","000000000000010011","000000000000001101","000000000000001111","000000000000001011","000000000000000011","000000000000001011","000000000000000000","111111111111110010","000000000001011000","111111111111011111","000000000000100110","111111111111100101","111111111111110000","000000000000001000","111111111111101111","000000000000000111","111111111111110010","111111111111101101","111111111111100000","111111111111110011","000000000000010100","000000000000011001","000000000000000100","000000000000010000","111111111111100101","000000000000101111","111111111111101011","000000000000001110","000000000000000100","111111111111111110","111111111111110101","000000000000100000","000000000000010001","000000000000000100","111111111111111000","111111111111111000","000000000000001000","000000000000100000","000000000000001010","000000000000010010","000000000000000110","111111111111101001","111111111111110000","000000000000011101","000000000000011100","111111111111100011","111111111111111101","000000000000100110","111111111111100110","000000000000001110","000000000000001001","000000000000010101","111111111111100110","000000000000010010","111111111111111010","000000000000010010","000000000000000000","000000000000010011","000000000000000101","000000000000001010","111111111111100010","111111111111100111","000000000000000000","000000000000100011","000000000000000110","000000000000001001","000000000000010100","111111111110111101","000000000000011011","111111111111110011","111111111111011100","000000000000000110","111111111111111001","111111111111110000","000000000000100011","000000000000001111","111111111111110010","000000000000000001","000000000000000111","000000000000010011","111111111111111000","111111111111110110","111111111110111101","111111111111111101","000000000000010101","000000000000011000","000000000000101000","000000000000000110","000000000000010001","000000000000101000","000000000000000101","000000000000001100","000000000000001101","000000000000001101","000000000000010001","000000000000100010","111111111111111110","111111111111110010","111111111111100111","000000000000000100","000000000000111101","000000000000001010","000000000000000110","111111111111100001","111111111111011011","000000000000010010","000000000000000000","111111111111111010","000000000000011101","111111111111101000","111111111111110111","000000000000000100","000000000000001010","111111111111111111","000000000000010000","000000000000000001","000000000000001000","000000000000000010","111111111111101101","111111111111100000","111111111111111101","111111111111111001","000000000000111010","000000000000000000","111111111111110000","111111111111101011","000000000000000100"),
("000000000000010000","111111111111000011","000000000000000111","111111111111110110","111111111111010011","111111111111111111","111111111111101101","000000000000011001","111111111111111100","000000000001010001","111111111111001000","000000000000010101","111111111111010111","111111111111110100","000000000000001001","111111111111011110","000000000000001000","111111111111010110","111111111111001100","111111111111100111","111111111111100001","000000000000010101","111111111111110100","000000000000000111","000000000000010001","000000000000000000","000000000000110000","111111111111100000","000000000000001011","000000000000010000","000000000000000101","111111111111110110","000000000000001101","000000000000000111","000000000000000000","000000000000100010","111111111111110100","111111111111100110","000000000000011100","111111111111111010","111111111111111010","111111111111101111","111111111111100100","000000000000001011","000000000000011111","000000000000110111","111111111111011011","000000000000100101","000000000000001101","111111111111110001","111111111111111101","000000000000001011","000000000000000011","111111111111101101","000000000000000110","111111111111101101","000000000000001000","111111111111101100","000000000000000101","111111111111111000","000000000000010011","111111111111110000","111111111111111010","111111111111100010","000000000000001100","000000000000000100","111111111111101011","000000000000011011","111111111110111101","000000000000011001","111111111111110101","111111111111011111","000000000000000111","111111111111111011","111111111111110010","000000000000100101","111111111111111100","111111111111110101","000000000000010111","000000000000000000","000000000000001000","000000000000010101","111111111111110000","111111111110100001","111111111111110111","000000000000101110","000000000000011010","000000000000011001","000000000000100110","000000000000000101","000000000000010110","000000000000000000","000000000000001101","000000000000000101","000000000000001100","111111111111101100","000000000000101010","111111111111110011","000000000000001101","111111111111101010","111111111111110111","000000000000101010","000000000000001000","111111111111111001","000000000000001101","111111111111101011","000000000000001101","000000000000001010","111111111111100010","000000000000011111","111111111111111101","111111111111101011","000000000000010101","000000000000011001","111111111111011110","000000000000001110","111111111111110000","000000000000010010","000000000000010110","111111111111110000","111111111111101001","000000000000010101","000000000000001110","000000000000101011","000000000000110011","000000000000000111","111111111111100110","000000000000001011"),
("000000000000011011","111111111110101100","000000000000000000","111111111111101111","111111111111100001","111111111111111000","000000000000000011","000000000000001101","111111111111101110","000000000000010010","111111111110111101","000000000000001000","111111111111011011","111111111111111101","111111111111111100","111111111111011111","000000000000100111","111111111111101011","111111111111101001","000000000000011011","111111111111111001","000000000000000100","111111111111110000","000000000000100110","000000000000011101","000000000000001010","000000000000110100","111111111111001011","000000000000001110","000000000000011100","111111111111101011","111111111111101100","000000000000000110","111111111111111100","000000000000001101","000000000000110001","111111111111111010","000000000000000110","000000000000001111","000000000000011110","000000000000000000","000000000000001001","111111111111111110","111111111111110100","000000000000001011","000000000000111110","000000000000000110","000000000000100110","000000000000100111","000000000000001111","000000000000100000","000000000000110101","000000000000000000","000000000000001000","000000000000001101","111111111111111011","000000000000001001","111111111111101110","000000000000001001","000000000000000101","111111111111101011","000000000000000111","000000000000000101","000000000000000000","000000000000110101","000000000000000110","111111111111110010","000000000000000000","111111111111001001","000000000000011010","111111111111101110","111111111111010001","111111111111111010","000000000000010001","111111111111111111","000000000000101000","000000000000010110","111111111111100010","111111111111111101","000000000000101001","000000000000101111","111111111111110001","000000000000001101","111111111110101001","000000000000000000","000000000000111111","000000000000100000","000000000000101001","000000000000010001","000000000000001100","000000000000011001","000000000000000101","111111111111110011","111111111111111111","111111111111111111","111111111111101110","000000000000101101","111111111111011111","000000000000100000","111111111111011011","111111111111010110","000000000000011110","111111111111101000","000000000000011001","000000000000011011","000000000000000111","111111111111101111","111111111111101010","000000000000000110","000000000000010101","111111111111110100","111111111111011111","000000000000001010","000000000000010000","111111111111111001","111111111111111100","000000000000010001","111111111111111000","000000000000100010","000000000000000010","111111111111011001","000000000000000000","000000000000000010","000000000000010101","000000000001000000","000000000000010111","111111111111000110","000000000000010001"),
("000000000000011100","111111111110110000","111111111111111101","111111111111101110","111111111111110111","111111111111101110","111111111111011010","111111111111110110","111111111111110101","111111111111100010","111111111111000111","111111111111101010","111111111111100010","000000000000000001","111111111111000010","111111111111110100","000000000000101110","111111111111101010","111111111111010101","111111111111101111","111111111111111110","111111111111110100","111111111111011010","000000000000101111","111111111111110100","111111111111111001","000000000000001101","111111111110111101","000000000000001000","000000000000010011","000000000000000011","111111111111110101","000000000000010010","111111111111110111","111111111111111001","000000000000010111","111111111111100101","000000000000011011","111111111111111110","111111111111111000","111111111111101011","000000000000100000","111111111111110001","000000000000000000","000000000000001010","000000000000001010","000000000000100011","000000000000011111","000000000000101010","000000000000100110","000000000000100100","000000000000001100","000000000000000000","000000000000000001","111111111111100011","111111111111101101","000000000000010011","111111111111101111","111111111111101011","111111111111111101","000000000000100011","111111111111110000","111111111111101110","111111111111111101","000000000000101000","000000000000000101","000000000000001110","111111111111111111","111111111111010011","111111111111111101","000000000000000011","111111111111011101","000000000000111001","111111111111110010","000000000000001101","000000000000110011","000000000000001100","111111111111101111","111111111111110000","000000000000000011","000000000000011100","000000000000001000","000000000000001001","111111111111010111","000000000000011010","000000000000010101","000000000000000101","000000000000100010","111111111111110100","000000000000101011","000000000000000001","000000000000010010","111111111111111011","000000000000000111","111111111111111011","000000000000001100","000000000000101100","111111111111110100","000000000000110001","111111111111111000","111111111111101010","000000000000000000","000000000000001000","000000000000101001","000000000000000110","000000000000010111","111111111111110100","111111111111000110","000000000000000100","111111111111100111","000000000000010111","111111111111010010","000000000000001000","000000000000001101","111111111111011001","111111111111100000","000000000000001001","111111111111111010","000000000000010100","000000000000000001","111111111111100100","000000000000001000","111111111111110100","111111111110110111","000000000000100000","111111111111111100","111111111111011010","000000000000011010"),
("111111111111111101","111111111111101011","111111111111111000","111111111111110111","000000000000010000","111111111111100010","111111111111101011","111111111111110110","000000000000011100","111111111111010011","111111111111010101","111111111111011011","111111111111110000","000000000000011100","111111111111100101","111111111111001111","000000000000001110","000000000000001100","111111111111100100","111111111111101011","000000000000101000","111111111111111011","111111111111001000","000000000000010011","000000000000000000","000000000000011111","111111111111011001","111111111111111011","000000000000010010","000000000000010101","000000000000010100","000000000000010110","111111111111101111","111111111111101001","000000000000001001","000000000000010101","111111111111110111","000000000000000011","111111111111110011","000000000000001100","111111111111111101","000000000000001111","000000000000011011","000000000000001010","000000000000000001","000000000000000000","000000000000101111","111111111111110110","111111111111110110","000000000000100110","000000000000100101","111111111111111001","111111111111011001","000000000000011010","000000000000000100","111111111111100010","000000000000010111","111111111111101011","000000000000000101","111111111111111101","000000000000110001","111111111111111101","111111111111010100","000000000000001011","000000000000101110","000000000000000001","000000000000010100","111111111111110101","000000000000000100","111111111111000100","000000000000101100","000000000000000000","000000000000011011","000000000000100111","000000000000100110","000000000000001111","111111111111100101","111111111111110001","111111111111110001","111111111111110001","000000000000000101","111111111111101110","111111111111101001","000000000000001011","000000000000001010","111111111111110110","111111111111111100","000000000000011111","111111111111010000","000000000000101111","000000000000000000","000000000000011111","111111111111111111","111111111111111011","111111111111111001","000000000000010110","000000000000010001","111111111111111000","000000000000001010","111111111111100001","111111111111011100","111111111111011100","000000000000011100","000000000000100110","000000000000011110","000000000000000110","000000000000010110","111111111111010001","000000000000010101","111111111111110100","000000000000001001","111111111111010101","000000000000000110","000000000000001100","111111111111111000","111111111111111010","000000000000001010","111111111111100110","111111111111111111","000000000000000000","111111111111110000","000000000000000001","000000000000011010","111111111110111101","000000000000101001","000000000000000010","111111111111100111","000000000000010011"),
("000000000000001010","111111111111110011","000000000000001000","000000000000001111","000000000000010010","111111111111101010","111111111111100011","000000000000000010","000000000000001000","111111111111100110","111111111111001111","111111111111011110","000000000000001001","000000000000010100","000000000000001100","111111111111011101","111111111111110101","111111111111110010","111111111111111100","111111111111010010","111111111111111010","000000000000010110","111111111111000101","000000000000011101","111111111111100110","111111111111111011","000000000000010000","000000000000001110","000000000000011010","111111111111110001","000000000000010000","000000000000001100","000000000000001001","111111111111111011","000000000000000111","000000000000001010","111111111111111100","000000000000010000","000000000000001001","111111111111110111","111111111111111000","000000000000001100","000000000000011010","000000000000100100","000000000000011000","111111111111111110","000000000000001001","111111111111111101","000000000000011111","000000000000100110","000000000000000000","111111111111111010","111111111111101101","000000000000001100","000000000000011000","111111111111111000","000000000000010110","111111111111101010","000000000000001000","111111111111111100","000000000000001010","000000000000000010","111111111111010010","111111111111110100","000000000000110001","111111111111111000","000000000000011111","111111111111110101","000000000000001000","111111111110111010","111111111111111111","111111111111101010","111111111111110111","000000000000010010","000000000000110110","111111111111110111","111111111111101011","111111111111101011","000000000000000110","111111111111111110","000000000000000000","111111111111101110","111111111111101100","000000000000100001","111111111111110111","111111111111110001","111111111111110100","111111111111111011","111111111111010011","000000000000001100","000000000000000010","111111111111111001","000000000000010110","111111111111100010","111111111111111100","000000000000101111","111111111111010110","111111111111110101","111111111111101111","000000000000000010","111111111111101100","111111111111011111","000000000000000011","111111111111111110","000000000000010100","111111111111111110","000000000000010110","111111111111111010","000000000000000100","111111111111111011","111111111111111100","111111111111011111","000000000000010100","000000000000000011","000000000000001011","111111111111100010","000000000000001000","111111111111010110","000000000000011100","111111111111110100","111111111111101010","111111111111101000","000000000000110100","111111111111000111","000000000000001000","000000000000000000","111111111111010101","000000000000101010"),
("111111111111101101","000000000000010001","111111111111111100","000000000000000000","000000000000101000","111111111111111110","111111111111100101","111111111111101011","000000000000100101","111111111111110110","111111111111010110","111111111111101000","000000000000001110","111111111111111011","000000000000100010","111111111111100010","000000000000001000","111111111111100011","111111111111111011","111111111111011001","111111111111111000","000000000000011110","111111111111110001","000000000000000001","111111111111100000","000000000000000100","111111111111101100","000000000000000001","000000000000011010","111111111111010100","000000000000000000","000000000000101100","111111111111101101","111111111111111000","000000000000010001","000000000000000101","111111111111110010","000000000000000000","111111111111111010","111111111111111100","111111111111101100","000000000000001101","000000000000011010","000000000000001100","111111111111110011","000000000000011100","111111111111111110","000000000000101011","111111111111111010","000000000000000001","000000000000000010","111111111111100100","000000000000001000","000000000000000110","000000000000011011","000000000000001011","000000000000010000","111111111111110100","000000000000010000","000000000000000101","000000000000010000","000000000000010010","111111111111110100","111111111111110110","000000000001000100","111111111111111110","000000000000000101","111111111111111010","111111111111111111","111111111111011000","000000000000010001","111111111111111001","111111111111110101","000000000000001001","000000000000101010","111111111111111001","111111111111101110","000000000000000010","000000000000011011","000000000000000110","111111111111101010","111111111111100111","111111111111111111","000000000000010100","000000000000000011","000000000000011010","000000000000000001","000000000000000000","111111111111100111","111111111111101000","000000000000001101","000000000000001100","000000000000101000","111111111111010110","000000000000010100","000000000000000011","111111111111011111","000000000000101011","111111111111011011","000000000000101001","111111111111101100","111111111111100000","111111111111110000","111111111111110100","111111111111101111","111111111111110000","111111111111111010","111111111111111001","000000000000010111","111111111111101100","111111111111111110","111111111111010100","000000000000010111","111111111111111110","000000000000001010","111111111111010101","000000000000000000","111111111111101101","000000000000000101","111111111111011100","111111111111111111","111111111111011111","000000000000110001","000000000000001001","000000000000001101","111111111111110101","111111111111100011","000000000000011001"),
("111111111111110100","000000000000010000","111111111111110100","111111111111101000","000000000000000001","111111111111101111","111111111111111110","111111111111111010","000000000000011010","000000000000001100","000000000000000111","111111111111101011","000000000000011000","111111111111111110","000000000000010010","111111111111101011","000000000000001001","111111111111111101","111111111111110100","111111111111101100","000000000000000001","000000000000001111","000000000000010001","111111111111110011","111111111111101001","111111111111111001","000000000000000011","000000000000001011","111111111111100110","111111111111011001","111111111111101101","000000000000011110","111111111111111000","000000000000010111","111111111111100000","000000000000001001","111111111111011001","111111111111110010","111111111111111011","111111111111110111","111111111111101100","000000000000000111","000000000000100110","000000000000100110","000000000000001110","111111111111111011","111111111111101110","111111111111111010","000000000000010000","000000000000000010","000000000000001011","111111111111101100","000000000000010101","000000000000000000","000000000000100011","111111111111110101","000000000000001001","111111111111101000","000000000000001110","000000000000001101","000000000000001101","111111111111111001","000000000000000101","000000000000001011","000000000000110100","000000000000001101","111111111111110010","111111111111111001","111111111111110110","000000000000010001","000000000000000000","111111111111101010","111111111111101101","000000000000100001","000000000000011110","000000000000000111","000000000000000001","000000000000001001","111111111111110110","000000000000000100","000000000000001100","000000000000010010","000000000000000100","000000000000000111","000000000000010010","000000000000001000","111111111111111101","000000000000001100","000000000000001011","111111111110111100","111111111111110100","000000000000000001","000000000000011010","111111111111010011","000000000000000001","000000000000001001","111111111111010001","000000000000100011","111111111111110001","000000000000111100","000000000000000000","111111111111101101","000000000000000011","000000000000010010","000000000000000001","111111111111101011","000000000000100100","111111111111111100","000000000000010000","000000000000000101","111111111111111000","111111111111101111","111111111111111011","000000000000011000","111111111111111000","111111111111110101","000000000000000111","111111111111110110","111111111111110011","111111111111110001","000000000000000010","111111111111111011","000000000000011111","000000000000100010","111111111111111100","000000000000001000","111111111111100011","000000000000001100"),
("111111111111101100","111111111111111011","000000000000000011","111111111111111111","111111111111010100","111111111111100110","111111111111111011","000000000000000010","111111111111110100","000000000000010001","000000000000010100","111111111111111000","111111111111110110","000000000000010011","000000000000000000","111111111111100110","000000000000000100","111111111111111010","111111111111100011","000000000000000111","111111111111111101","000000000000000000","000000000000001110","111111111111100101","000000000000000101","111111111111110000","111111111111111111","000000000000011110","111111111111111100","111111111111101111","111111111111110110","000000000000100101","000000000000010000","000000000000001000","111111111111100110","000000000000011100","111111111111100101","111111111111110100","111111111111100011","000000000000011100","000000000000001100","000000000000000101","000000000000010000","000000000000011100","000000000000010001","111111111111110111","000000000000000010","000000000000010011","111111111111110111","000000000000000111","111111111111101000","000000000000001000","111111111111111100","000000000000010010","000000000000011001","111111111111110111","000000000000010001","000000000000010100","000000000000011001","000000000000001111","000000000000010000","000000000000001010","111111111111110110","000000000000001010","000000000000000001","000000000000010011","111111111111111011","111111111111101111","111111111111110111","000000000000001010","111111111111110111","111111111111101010","111111111111110111","000000000000101101","000000000000000011","000000000000001000","000000000000001010","000000000000000100","000000000000010000","111111111111101101","111111111111101110","000000000000001101","111111111111111010","000000000000000111","000000000000000100","000000000000110011","000000000000011110","111111111111110110","000000000000000011","111111111111010011","000000000000000100","111111111111101101","000000000000011001","111111111111110010","000000000000010111","000000000000001001","111111111111001000","111111111111111111","000000000000011001","000000000000110111","111111111111100000","000000000000000011","111111111111101010","000000000000001110","000000000000010000","111111111111110101","000000000000000001","111111111111111101","000000000000001001","000000000000001001","000000000000010010","111111111111101001","111111111111111011","000000000000001011","000000000000010100","111111111111111011","111111111111111101","000000000000011001","000000000000000000","000000000000000110","111111111111110001","111111111111100010","111111111111111100","000000000000001011","000000000000010111","000000000000011011","111111111111111111","000000000000011011"),
("111111111111010011","000000000000000100","111111111111110111","000000000000001101","111111111111001010","111111111111110011","000000000000001010","111111111111111101","000000000000000000","000000000000000000","000000000000001010","111111111111111001","000000000000001111","000000000000101011","111111111111111110","111111111111100001","111111111111100100","111111111111110111","111111111111100100","111111111111110000","000000000000000010","111111111111111001","111111111111101111","111111111111110110","000000000000000110","000000000000000110","111111111111110111","000000000000001100","111111111111110001","111111111111001110","111111111111111111","000000000000011110","000000000000101010","111111111111111111","111111111111001001","000000000000011000","111111111111110011","000000000000010011","000000000000000000","111111111111110010","000000000000000000","000000000000001110","000000000000000111","000000000000110100","000000000000011010","111111111111011001","000000000000011001","000000000000000110","111111111111110110","111111111111101011","111111111111111101","000000000000100101","000000000000000000","000000000000001101","111111111111111101","000000000000000001","111111111111101100","000000000000010001","000000000000001010","000000000000000000","000000000000000000","111111111111101000","000000000000001111","000000000000100001","111111111111100101","111111111111111111","111111111111110001","000000000000001100","000000000000000011","000000000000001011","111111111111110111","111111111111110101","111111111111101000","000000000000000001","000000000000010000","111111111111101010","000000000000001111","000000000000001011","000000000000010011","000000000000001111","111111111111101010","000000000000010101","000000000000000100","111111111111101010","000000000000010000","000000000000011011","000000000000100010","111111111111011110","000000000000000110","111111111111101011","111111111111111000","000000000000000101","000000000000000011","000000000000000101","000000000000010010","111111111111111010","111111111111010111","000000000000000110","111111111111110000","000000000000101111","000000000000001110","000000000000010000","111111111111111100","000000000000010100","111111111111110011","000000000000001011","000000000000001110","000000000000010110","000000000000001100","000000000000000011","000000000000001101","111111111111111011","000000000000000111","000000000000000000","000000000000100101","000000000000000101","000000000000000000","111111111111110011","111111111111111110","000000000000001000","111111111111001111","111111111111101101","111111111111110000","111111111111111111","000000000000001000","111111111111110101","111111111111010111","111111111111110111"),
("111111111111000010","000000000000000111","000000000000000001","000000000000010001","111111111111100011","000000000000000010","000000000000000001","111111111111110011","111111111111110101","111111111111110111","111111111111101100","000000000000000000","111111111111110000","000000000000000000","000000000000010001","000000000000000000","111111111111110000","111111111111110100","111111111111101011","111111111111110111","111111111111110000","000000000000001101","111111111111110010","000000000000001100","111111111111110101","111111111111111000","111111111111111010","000000000000100011","111111111111110111","111111111111010100","111111111111110010","000000000000001111","000000000000000111","111111111111110110","111111111111111101","000000000000000000","111111111111011110","111111111111111001","000000000000010001","111111111111100111","000000000000001010","000000000000110100","111111111111110011","000000000000001000","000000000000010110","111111111111110000","000000000000100111","111111111111110011","000000000000001101","111111111111111011","000000000000000010","000000000000001001","111111111111110111","000000000000001100","111111111111111001","000000000000010000","111111111111101011","000000000000010101","000000000000000010","111111111111101111","000000000000001111","000000000000001001","000000000000010111","111111111111111101","111111111111011100","000000000000011101","111111111111100111","111111111111101111","111111111111011111","111111111111111110","000000000000010001","111111111111101101","111111111111011110","111111111111100011","000000000000001101","111111111111100011","000000000000001001","000000000000010010","000000000000010000","111111111111110111","000000000000001110","000000000000011011","111111111111101111","000000000000000111","000000000000010000","000000000000001110","000000000000111001","111111111111010100","000000000000010110","111111111111110110","111111111111100110","000000000000000010","111111111111111100","000000000000000110","000000000000001110","111111111111110101","111111111111100101","000000000000000001","111111111111111011","000000000000110111","000000000000001101","000000000000000011","111111111111101001","000000000000000100","111111111111110110","000000000000011010","000000000000000101","000000000000001100","000000000000011111","111111111111110110","000000000000010011","000000000000100010","111111111111111011","000000000000011000","000000000000001101","000000000000010100","000000000000001101","111111111111111010","000000000000011011","111111111111110101","111111111111001111","111111111111111101","111111111111010111","000000000000001111","000000000000000100","111111111111110101","111111111111101010","111111111111110000"),
("111111111111010100","111111111111111001","111111111111111110","000000000000011110","000000000000000100","000000000000000010","000000000000101000","111111111111100000","111111111111111010","111111111111100101","111111111111101010","111111111111100010","111111111111011101","111111111111101100","000000000000100110","111111111111111001","000000000000000010","111111111111110011","111111111111111110","111111111111011101","000000000000010001","000000000000111010","000000000000000100","000000000000101000","111111111111110011","000000000000010000","000000000000011000","111111111111101111","111111111111110001","111111111111011111","111111111111101100","000000000000101101","000000000000000111","111111111111100001","111111111111111101","111111111111101111","111111111111010111","111111111111010001","111111111111110110","111111111111100010","111111111111110000","000000000000001010","000000000000001011","000000000000000010","000000000000000000","111111111111101010","000000000000001001","000000000000100100","111111111111111011","000000000000010110","000000000000000000","111111111111111011","000000000000000110","111111111111110101","111111111111010110","000000000000011101","111111111111100001","000000000000001010","111111111111111100","111111111111110101","000000000000001011","111111111111111001","000000000000001010","000000000000000110","111111111111001110","111111111111111000","111111111111011110","000000000000010010","111111111111011110","111111111111100100","000000000000011111","111111111111110001","111111111111100110","111111111111100001","111111111111110010","111111111111110110","000000000000000001","000000000000001111","000000000000001111","000000000000010010","000000000000000110","000000000000010011","111111111111101010","000000000000011000","000000000000000101","111111111111111011","000000000000110000","111111111111001111","000000000000000001","111111111111111000","000000000000001010","111111111111110000","000000000000001000","000000000000010001","000000000000010100","111111111111101111","000000000000001010","111111111111110010","111111111111001111","000000000000000101","000000000000001000","000000000000100000","000000000000000111","000000000000000001","000000000000010011","000000000000011011","111111111111110111","000000000000101010","000000000000010101","111111111111110010","111111111111111101","000000000000011011","111111111111111000","111111111111101001","000000000000010001","000000000000100100","111111111111111001","111111111111100101","000000000000000101","111111111111101100","111111111110110100","000000000000001111","111111111111110000","000000000000000111","000000000000010101","000000000000000100","111111111111010111","111111111111111110"),
("111111111110100110","111111111111111111","111111111111110111","111111111111111110","111111111111101101","111111111111110101","000000000000011001","111111111111100001","111111111111110000","000000000000100000","111111111111110001","111111111111101011","111111111111011110","111111111111000101","000000000000001001","111111111111111101","000000000000001000","000000000000000001","111111111111101001","111111111111110000","000000000000010110","000000000000110000","000000000000010101","000000000000010111","000000000000000000","000000000000000101","000000000000000110","000000000000000011","000000000000000100","111111111111101001","111111111111011100","000000000000110110","111111111111111101","111111111111011000","000000000000000001","111111111111010101","111111111111000011","111111111111100000","000000000000000000","111111111111011100","111111111111111011","000000000000001001","111111111111111110","111111111111010000","111111111111011011","111111111111100110","000000000000001100","000000000000000001","111111111111111111","000000000000100101","000000000000010101","111111111111100100","000000000000010111","000000000000010101","111111111111111011","111111111111110010","111111111111001111","111111111111110101","000000000000011100","000000000000001001","000000000000010011","111111111111111011","111111111111101111","000000000000000111","111111111111011000","000000000000001010","111111111111110110","111111111111111111","111111111111101110","111111111111111101","111111111111110010","111111111111100110","111111111111101000","111111111111001100","000000000000010010","000000000000000100","000000000000000000","000000000000000001","000000000000011110","000000000000001000","000000000000000110","111111111111100011","000000000000000001","111111111111101010","111111111111111011","111111111111110110","000000000000101000","111111111111010001","111111111111110100","000000000000000011","111111111111111101","000000000000000100","000000000000100001","000000000000100000","000000000000000001","000000000000000011","111111111111110110","000000000000000111","111111111111010000","111111111111110111","000000000000010010","000000000000011000","000000000000100000","111111111111110101","000000000000001110","000000000000001111","000000000000001100","000000000000100100","000000000000011011","000000000000010111","000000000000000110","000000000000011101","000000000000001010","111111111111100111","000000000000011010","000000000000100110","000000000000000101","111111111111100001","000000000000000100","111111111111100000","111111111111000011","000000000000001101","111111111111011101","000000000000011001","000000000000010110","111111111111101101","111111111111011100","111111111111111110"),
("111111111110100010","000000000000110000","111111111111101110","111111111111111010","000000000000000011","000000000000001011","000000000000100101","000000000000010001","111111111111111010","000000000000010100","111111111111010000","111111111111111011","111111111111100111","111111111111000110","111111111111111111","111111111111110001","111111111111110101","111111111111110001","000000000000001001","111111111111110101","000000000000101010","000000000000010101","000000000000000110","000000000000101111","000000000000001110","111111111111110011","111111111111011111","000000000000000000","000000000000001100","111111111111111100","111111111111001011","000000000000011111","000000000000000010","111111111111101000","111111111111111011","111111111111100111","111111111110110100","111111111111010010","000000000000011011","111111111110111000","000000000000000111","000000000000000000","111111111111101010","111111111111011110","111111111111100100","000000000000000000","111111111111110111","000000000000000111","111111111111110011","000000000000011000","111111111111111101","111111111111011101","000000000000100001","000000000000001101","111111111111100101","000000000000001111","111111111111100101","000000000000000101","000000000000001011","111111111111111110","000000000000010010","111111111111011101","111111111111001101","000000000000000001","111111111111001100","000000000000100001","111111111111111110","000000000000010011","000000000000001100","111111111111101001","000000000000001110","111111111111001001","111111111111100110","111111111111011010","000000000000011000","111111111111110110","000000000000000001","111111111111101101","111111111111111011","000000000000000111","000000000000011010","000000000000000010","111111111111110111","111111111111101101","111111111111100101","111111111111011110","000000000000000000","111111111111010111","111111111111110010","000000000000100100","111111111111110110","000000000000011110","000000000000111000","000000000000011010","000000000000010000","111111111111110010","111111111111111001","000000000000011001","111111111111000000","111111111111001111","000000000000001110","000000000000110000","000000000000100100","111111111111101111","000000000000010001","000000000000101001","000000000000011010","000000000000011101","000000000000001110","111111111111101010","000000000000010111","000000000000101100","000000000000001111","111111111111001001","000000000000000101","000000000000010010","000000000000100100","111111111111100100","000000000000100101","111111111111111000","111111111110101111","111111111111111111","111111111111010000","111111111111010111","111111111111111000","000000000000010110","111111111111000110","000000000000001001"),
("111111111110110111","000000000000011100","111111111111011111","111111111111101001","111111111111110010","111111111111111111","000000000000010111","000000000000001010","000000000000001000","000000000000100000","000000000000011010","000000000000011101","111111111111111110","111111111111101001","111111111111101110","000000000000000001","111111111111111100","000000000000011001","111111111111111101","000000000000001101","111111111111101101","111111111111110101","000000000000010000","000000000000001010","000000000000001010","000000000000001110","000000000000011111","111111111111111001","000000000000100011","000000000000000010","111111111111100001","000000000000001110","111111111111111100","111111111111101000","000000000000001011","111111111111110010","111111111111000001","111111111111011101","111111111111111111","111111111110100111","111111111111101110","000000000000000001","111111111111010111","111111111111011011","111111111111101100","111111111111111010","000000000000101000","000000000000100101","111111111111010011","111111111111011100","000000000000101100","111111111111101101","000000000000010101","111111111111000011","111111111111010010","111111111111100101","111111111111010110","111111111111111101","111111111111101100","000000000000010101","111111111111101000","000000000000000110","111111111111100010","000000000000000011","111111111111010101","000000000000000000","111111111111110111","000000000000100110","000000000000000101","111111111111101111","000000000000011110","111111111111100000","000000000000000010","111111111111101110","111111111111100110","000000000000000111","000000000000010100","111111111111011100","111111111111100010","000000000000110011","000000000000000010","111111111111011001","111111111111111101","111111111111110000","111111111111110101","111111111111011000","111111111111001110","111111111111011000","111111111111010101","111111111111011100","111111111111001110","000000000000001101","000000000000011001","000000000000000100","111111111111001110","111111111111001000","111111111111111111","000000000000100111","111111111110101110","111111111111010111","000000000000011000","000000000000101111","111111111111101101","000000000000001011","000000000000010011","000000000000101111","111111111111100000","111111111111110000","000000000000000010","111111111111100011","111111111111110100","000000000000010010","000000000000010011","111111111111010010","111111111111101000","000000000000101001","000000000000111011","111111111111011111","000000000000100110","111111111111001110","111111111110100010","000000000000001001","111111111111110100","111111111111110010","000000000000001001","000000000000001000","000000000000001100","111111111111101110"),
("111111111111000110","111111111111100110","000000000000001001","111111111111111010","000000000000000000","111111111111101101","111111111111110101","000000000000001010","000000000000011100","111111111111101111","000000000000100000","000000000000011110","111111111111111001","000000000000001010","111111111111100111","000000000000000100","111111111111101011","000000000000011010","000000000000011011","111111111111111100","000000000000010000","111111111111100111","111111111111100000","111111111111010111","111111111111110110","000000000000000011","000000000000000101","111111111111100111","000000000000001000","111111111111111000","111111111111111011","000000000000010101","111111111111110001","111111111111100101","000000000000110101","111111111111110100","111111111111101111","000000000000001100","000000000000001010","111111111111011100","111111111111011110","000000000000000100","111111111111110011","111111111111011010","111111111111101010","111111111111111101","000000000000010100","000000000000011100","000000000000001110","111111111111101101","000000000000010100","000000000000001111","111111111111101001","111111111111101000","000000000000001000","000000000000001011","111111111111110101","111111111111110000","111111111111011100","111111111111101111","111111111111101100","111111111111110100","000000000000001001","111111111110111101","111111111111101011","111111111111101110","000000000000110010","000000000000001111","000000000000011010","111111111111111110","111111111111111100","000000000000001101","000000000000001011","000000000000000010","111111111111011100","000000000000000011","000000000000010110","111111111111100001","111111111111101101","000000000000010010","111111111111100011","000000000000000110","111111111111110000","000000000000001001","000000000000000010","111111111111110000","111111111111110100","111111111111010001","111111111111000000","111111111111100111","111111111111000111","111111111111100001","000000000000101101","111111111111101011","111111111111011110","111111111111011110","000000000000011001","000000000000010100","111111111111101001","111111111111001010","000000000000010110","111111111111111000","111111111111010110","111111111111110100","000000000000100101","000000000000011011","111111111111110110","111111111111101011","111111111111111001","111111111111000110","111111111111101001","111111111111101111","111111111111101011","000000000000000100","000000000000000110","111111111111100011","000000000000001001","000000000000001011","111111111111111000","111111111111110001","111111111111011100","000000000000000101","000000000000001011","111111111111111001","111111111111110101","111111111111100001","111111111111111111","111111111111111011"),
("111111111111100011","111111111111101001","000000000000101010","111111111111101000","111111111111101111","111111111111010000","111111111111011011","111111111111011110","000000000000000000","111111111111100110","000000000000100110","000000000000010010","111111111111111010","000000000000000001","111111111111100110","000000000000001001","111111111111011010","000000000000010011","111111111111110000","000000000000000110","000000000001000000","111111111111111111","111111111111101010","000000000000000100","000000000000100000","000000000000000111","111111111111111111","111111111111101110","111111111111111111","000000000000000111","000000000000011001","111111111111100111","000000000000011010","000000000000000111","000000000000101011","111111111111101001","111111111111111000","000000000000100111","111111111111100000","000000000000010100","111111111111111100","000000000000011100","000000000000001011","111111111111011001","000000000000000010","111111111111100111","000000000000001010","000000000000010011","000000000000100010","111111111111100101","111111111111110101","000000000000010100","111111111111110101","000000000000101000","000000000000100101","000000000000011110","111111111111110101","111111111111111111","111111111111100010","000000000000000011","000000000000011101","000000000000010000","111111111111110011","111111111111010101","111111111111000011","000000000000001011","000000000000111011","111111111111011111","000000000000000001","000000000000011011","111111111111110101","111111111111101111","000000000000111000","111111111111101101","111111111111110001","111111111111110001","000000000000010100","111111111111111011","111111111111001001","111111111111111000","111111111111011110","000000000000001111","111111111111011100","111111111111110111","000000000000001110","111111111111100110","000000000000010111","111111111111110101","111111111111011011","000000000000000000","111111111111100001","111111111111100010","000000000000110011","111111111111010011","111111111111110110","111111111111100110","111111111111101110","000000000000011011","000000000000000101","111111111111110000","000000000000000000","111111111111111011","111111111111010100","000000000000000001","000000000000011010","111111111111111001","111111111111110111","111111111111100001","111111111111101111","111111111111101010","111111111111111101","111111111111111101","111111111111011001","111111111111100101","000000000000001101","111111111111011101","111111111111011000","000000000000001000","000000000000010011","111111111111110100","111111111111111000","111111111111111011","000000000000000000","111111111111011110","111111111111111100","111111111111011000","111111111111110010","111111111111111101"),
("111111111111010001","000000000000000000","111111111111111111","000000000000000100","111111111111100100","111111111111101010","000000000000100101","111111111111111000","000000000000001111","000000000000000011","111111111111111100","111111111111111000","000000000000000110","000000000000011010","000000000000000100","000000000000000011","111111111111111001","000000000000000100","000000000000000000","111111111111111110","000000000000100000","111111111111110111","111111111111101001","111111111111110101","111111111111111101","111111111111100111","111111111111010000","111111111111111100","000000000000001011","111111111111111011","000000000000000100","000000000000000011","111111111111110010","111111111111110000","000000000000011111","111111111111111011","000000000000000111","000000000000001100","111111111111011110","000000000000000111","111111111111110000","000000000000000000","000000000000101100","111111111111101100","111111111111110100","000000000000010001","000000000000010100","111111111111111010","000000000000001101","000000000000010101","000000000000000001","111111111111100111","000000000000000011","000000000000100101","000000000000000010","000000000000001101","111111111111111100","111111111111111111","000000000000010001","000000000000001010","111111111111111011","000000000000000100","000000000000000001","111111111111110000","000000000000000001","000000000000010000","111111111111100111","111111111111010010","111111111111110010","111111111111110010","111111111111101011","111111111111111010","000000000000100001","111111111111101011","111111111111111110","111111111111111100","111111111111110000","111111111111100110","000000000000010111","111111111111101001","111111111111011001","111111111111101110","111111111111110110","000000000000110000","111111111111110011","000000000000011011","000000000000000111","111111111111101010","111111111111101010","000000000000101010","111111111111111110","111111111111101100","000000000000010011","111111111111110001","000000000000011010","111111111111010101","000000000000001000","000000000000011100","111111111111110000","000000000000100110","111111111111100000","111111111111110001","111111111111100101","111111111111101111","000000000000011100","111111111111111010","111111111111110000","000000000000011000","111111111111111000","000000000000011001","000000000000001011","111111111111110011","111111111111010010","111111111111110100","000000000000010001","000000000000000111","111111111111011010","000000000000001010","111111111111010101","111111111111110010","111111111111101011","111111111111101100","000000000000011010","111111111111110110","000000000000010011","111111111111111100","000000000000000010","000000000000000100"),
("000000000000000001","111111111111110101","111111111111110001","000000000000001100","111111111111111010","000000000000000010","000000000000000111","111111111111111100","000000000000000000","000000000000001100","000000000000011001","111111111111111110","111111111111110010","000000000000010010","111111111111101101","000000000000001100","111111111111110110","111111111111110100","000000000000001000","000000000000000010","000000000000001101","000000000000001111","000000000000000011","000000000000010010","000000000000001111","111111111111111110","111111111111110100","111111111111111001","000000000000000010","000000000000011010","000000000000000000","111111111111111100","111111111111110111","111111111111111010","111111111111110011","111111111111111010","111111111111111000","000000000000000110","111111111111111111","111111111111110111","111111111111111001","000000000000001000","000000000000000100","000000000000000100","111111111111101001","000000000000000001","111111111111110100","000000000000001010","000000000000000110","111111111111111110","111111111111101111","111111111111101101","000000000000000010","000000000000000100","000000000000010000","111111111111111000","000000000000001010","111111111111111110","111111111111111001","111111111111110110","111111111111101001","000000000000001000","111111111111101100","000000000000001111","000000000000011101","000000000000001001","111111111111110011","000000000000001001","111111111111101000","111111111111111101","000000000000010111","000000000000001100","111111111111111001","111111111111111100","000000000000001010","000000000000000010","111111111111111101","000000000000000110","111111111111111101","111111111111101001","111111111111110110","111111111111101110","111111111111111110","000000000000000101","000000000000000011","000000000000001111","000000000000000000","000000000000001110","000000000000001011","000000000000011010","000000000000010000","111111111111110000","000000000000000010","000000000000010101","111111111111111000","111111111111110010","111111111111110110","111111111111101100","000000000000000101","111111111111111100","000000000000001111","000000000000001111","111111111111101010","000000000000001001","111111111111110110","000000000000010001","000000000000001000","111111111111110001","111111111111101111","000000000000001110","111111111111101011","111111111111111101","111111111111110110","111111111111101100","111111111111101101","111111111111111011","111111111111111100","111111111111110011","000000000000001000","111111111111111001","111111111111111001","111111111111110001","111111111111111000","111111111111101100","000000000000010011","000000000000010000","000000000000000001","111111111111111010"),
("000000000000001100","111111111111110010","111111111111111000","111111111111101010","111111111111111010","111111111111110000","111111111111110001","111111111111101100","111111111111111110","000000000000000100","000000000000100100","000000000000000000","000000000000001100","111111111111111011","000000000000010010","000000000000010111","111111111111111110","111111111111111001","111111111111110111","111111111111111010","000000000000100001","000000000000011000","000000000000011101","000000000000000000","000000000000010010","111111111111101010","111111111111110111","111111111111101111","000000000000010000","000000000000011000","000000000000000111","000000000000010100","000000000000000000","111111111111101100","000000000000010100","111111111111110010","000000000000011000","111111111111101110","111111111111101100","000000000000000110","000000000000011110","111111111111111111","000000000000010100","111111111111101111","111111111111100000","000000000000010001","111111111111111100","000000000000010001","000000000000000110","111111111111110111","000000000000000000","111111111111101000","000000000000100111","000000000000001000","000000000000001110","000000000000010111","111111111111110111","000000000000011000","000000000000000111","111111111111111101","111111111111110111","111111111111111001","111111111111111001","111111111111101001","111111111111110110","000000000000010000","000000000000000000","111111111111101000","000000000000010100","000000000000100001","111111111111011010","111111111111111100","000000000000010111","000000000000001010","111111111111101010","111111111111110000","000000000000000001","111111111111110111","000000000000000011","000000000000000101","000000000000001001","111111111111101110","111111111111100110","000000000000001001","111111111111110111","000000000000100011","000000000000000011","111111111111100001","000000000000000110","000000000000010110","000000000000010010","111111111111101110","000000000000010001","000000000000001000","000000000000010000","111111111111100101","111111111111111100","111111111111111001","000000000000001001","000000000000101000","000000000000010100","000000000000001001","111111111111111100","111111111111110110","000000000000001000","000000000000010101","111111111111110000","000000000000000011","000000000000000110","000000000000010001","111111111111111000","111111111111111010","111111111111110111","000000000000011101","111111111111111010","111111111111100101","111111111111100011","111111111111111111","111111111111110000","000000000000001110","000000000000010111","000000000000010100","111111111111100110","000000000000100001","000000000000000000","000000000000000100","000000000000001100","111111111111011110"),
("000000000000000111","111111111111101111","000000000000001110","111111111111011001","000000000000000100","111111111111011001","000000000000000001","111111111111011000","000000000000001000","000000000000011111","000000000000101100","000000000000001010","000000000000100010","000000000000000111","000000000000001100","000000000000000011","000000000000000011","000000000000010011","000000000000011111","000000000000000010","000000000000010100","000000000000011110","111111111111111000","111111111111111011","000000000000010111","111111111111011011","111111111111101110","111111111111011110","000000000000001100","111111111111111110","111111111111010100","000000000000001000","111111111111010101","111111111111101010","000000000000100010","111111111111110011","000000000000010011","111111111111101100","111111111111111011","000000000000000100","000000000000010100","000000000000101111","000000000000101001","111111111111101100","111111111111100110","000000000000001101","111111111111111110","111111111111101001","000000000000100001","000000000000001100","000000000000010010","111111111111011110","000000000000011000","111111111111110001","000000000000011110","000000000000001011","111111111111110011","111111111111111110","000000000000011110","111111111111111001","000000000000001010","111111111111111111","111111111111110111","111111111111011110","111111111111011000","000000000000010111","111111111111101110","111111111111111100","000000000000001011","000000000000100001","111111111111010010","111111111111110111","000000000000001001","000000000000101011","111111111111110110","111111111111101001","111111111111010100","111111111111110111","000000000000100001","000000000000000000","111111111111111010","111111111111011110","000000000000000101","000000000000100000","111111111111110111","000000000000100100","000000000000000111","111111111111100010","111111111111101001","000000000000010001","111111111111111100","111111111111100001","000000000000000111","000000000000000100","000000000000010010","111111111111100000","111111111111100010","111111111111101001","000000000000001000","000000000000110100","111111111111110001","111111111111111110","111111111111110001","111111111111110110","000000000000000111","111111111111101011","111111111111110100","111111111111111101","111111111111101010","000000000000001001","000000000000001110","000000000000000100","111111111111110011","000000000000010110","000000000000000110","111111111111101111","111111111111011011","000000000000000011","111111111111101100","000000000000001111","111111111111111111","000000000000000110","000000000000001101","000000000000100110","000000000000000100","111111111111101110","000000000000001000","111111111111010110"),
("000000000000001001","000000000000001000","000000000000000010","000000000000100001","000000000000010011","111111111111111010","111111111111111000","000000000000010111","000000000000001011","000000000000001011","111111111111011011","000000000000011001","000000000000001100","000000000000010111","000000000000001000","111111111111111110","111111111111011001","000000000000011100","111111111111100001","111111111111100111","111111111111110100","000000000000001011","000000000000000000","111111111111011101","000000000000001000","111111111111111111","111111111111101110","000000000000001010","111111111111111110","000000000000010011","000000000000000010","000000000000100000","111111111111110111","111111111111101010","111111111111111110","111111111111101000","111111111111100011","000000000000001111","111111111111101110","000000000000000011","111111111111111010","000000000000001101","000000000000100111","111111111111111101","111111111111111000","000000000000011001","000000000000000101","000000000000000000","000000000000001101","111111111111111011","111111111111111111","000000000000001010","000000000000011101","000000000000001110","000000000000010101","000000000000010001","111111111111111001","111111111111011000","000000000000011101","000000000000001001","000000000000000001","111111111111011101","111111111111110101","111111111111011110","000000000000001100","111111111111110011","000000000000011010","111111111111010000","111111111110111101","000000000000000000","111111111111111110","111111111111111000","000000000000000001","000000000000100001","111111111111100110","111111111111011111","111111111111101001","000000000000000010","111111111111110010","111111111111100010","111111111111011010","000000000000000100","111111111111110001","000000000000000001","000000000000011001","111111111111111100","000000000000000100","111111111111100011","111111111111011011","000000000000100000","111111111111100011","111111111111101000","000000000000100001","111111111111111111","000000000000100010","111111111111100001","111111111111101110","111111111111111001","000000000000001011","000000000000011100","111111111111100000","111111111111100110","111111111111111000","000000000000000000","000000000000000100","000000000000001010","000000000000001101","000000000000010011","111111111111101001","000000000000000100","000000000000010101","000000000000100011","111111111111110000","111111111111111111","000000000000001111","111111111111111110","000000000000000000","111111111111111010","111111111111011110","000000000000001011","111111111111100110","000000000000010100","000000000000011110","000000000000110001","111111111111110000","111111111111111111","111111111111101010","000000000000001000"),
("000000000000000011","000000000000011101","000000000000011111","000000000000000001","111111111111110010","111111111111011101","000000000000000101","000000000000010000","111111111111001101","111111111111111010","000000000000001001","000000000000000111","111111111111010011","000000000000001011","000000000000000101","111111111111011100","111111111111110000","111111111111101111","111111111111010101","111111111111011100","111111111111110011","000000000000101001","000000000000010100","111111111111011110","000000000000101001","000000000000000011","111111111111110111","111111111111100001","111111111111110010","000000000000000011","111111111111110101","000000000000010110","111111111111111100","000000000000000000","111111111111101110","111111111111111101","111111111111110100","111111111111110011","111111111111101101","111111111111100111","000000000000010111","000000000000100100","000000000000011110","111111111111101011","111111111111110000","111111111111110011","111111111111101000","111111111111011010","000000000000001111","000000000000000000","111111111111010100","111111111111100010","111111111111110110","111111111111111011","111111111111100011","000000000000011010","111111111111110100","111111111111010001","000000000000011000","111111111111110010","000000000000010000","111111111110111100","111111111111001110","000000000000000010","111111111111111100","000000000000001101","000000000000011000","111111111111100010","111111111110110100","111111111111010100","000000000000000100","111111111111101111","000000000000000100","000000000000011111","111111111111110101","111111111111011101","111111111111101011","000000000000000000","000000000000001010","111111111111100010","111111111111110010","000000000000011011","111111111111111100","111111111111110110","111111111111111011","111111111111011101","000000000000001100","111111111111101011","111111111111011100","111111111111110100","111111111111110000","000000000000010110","000000000000010100","111111111111110010","000000000000100111","000000000000000011","111111111111100010","111111111111111010","111111111111101110","000000000000110110","000000000000001001","111111111111110010","000000000000100010","000000000000001100","111111111111101111","111111111111111001","000000000000101110","000000000000000000","000000000000011110","111111111111111111","000000000000011111","000000000000101000","111111111111111111","111111111111101010","111111111111100001","000000000000010000","111111111111111001","111111111111110101","111111111111010011","111111111111011110","111111111111011101","111111111111101101","000000000000100110","111111111111111010","111111111111110000","111111111111100000","111111111111010001","000000000000011001"),
("000000000000000100","000000000000011101","000000000000100000","111111111111111010","000000000000010110","111111111111110111","000000000000000100","000000000000100100","111111111111001100","000000000000001011","000000000000001111","000000000000011001","111111111111011110","111111111111100001","000000000000001001","111111111111001001","000000000000000100","111111111111110000","111111111111001001","111111111111001111","000000000000000011","111111111111110111","000000000000000101","111111111111110001","000000000000010010","111111111111111110","000000000000001111","111111111111101011","111111111111111001","000000000000011000","000000000000000001","000000000000001001","000000000000001001","111111111111011011","111111111111110100","111111111111100111","111111111111111100","111111111111011100","111111111111111100","000000000000001000","111111111111111001","000000000000000000","000000000000000011","111111111111110000","111111111111111000","111111111111111100","000000000000000110","111111111111111111","000000000000010101","000000000000010011","111111111111011001","111111111111111110","000000000000010010","000000000000001100","111111111111100100","000000000000010011","111111111111011100","111111111111101001","000000000000100101","111111111111111110","000000000000010100","111111111111100000","111111111111010001","111111111111111100","111111111110101011","000000000000100010","000000000000000100","111111111111111111","111111111110010001","111111111111110111","000000000000001110","111111111111100100","000000000000011011","111111111111101010","000000000000010100","111111111111110010","000000000000001110","111111111111110110","111111111111110111","000000000000000011","000000000000000010","000000000000000001","111111111111110011","111111111111101011","111111111111101100","111111111111110011","000000000001000000","111111111111110110","111111111111001101","000000000000000111","111111111111011100","000000000000010010","000000000000010100","111111111111110011","000000000000011101","111111111111101110","000000000000001011","000000000000000100","111111111111110011","000000000000000011","000000000000011011","000000000000010100","111111111111110000","000000000000001100","111111111111100000","000000000000010001","000000000000000010","111111111111111111","111111111111100101","111111111111110100","000000000000001010","000000000000011001","000000000000001101","111111111111110001","000000000000000001","000000000000000000","111111111111111000","111111111111111000","111111111111010011","111111111111100101","111111111111010100","111111111111101101","111111111111111001","000000000000010101","111111111111100111","111111111111100101","111111111111010000","000000000000000010"),
("000000000000100101","000000000000011010","000000000000101001","000000000000001000","000000000000011001","000000000000001111","000000000000011101","000000000000001010","111111111111000100","000000000000111111","111111111111101101","000000000000101101","111111111111100101","000000000000000000","000000000000001111","111111111111010111","000000000000001100","000000000000000011","111111111111110101","111111111111100001","111111111111110100","000000000000011011","000000000000101001","111111111111111101","000000000000010011","000000000000000101","000000000000001011","000000000000000001","111111111111101111","111111111111110110","111111111111100010","000000000000001000","111111111111110001","111111111111010100","111111111111111011","000000000000010100","111111111111110111","111111111111101011","111111111111101001","111111111111101101","000000000000000101","111111111111100010","111111111111111001","111111111111011110","000000000000010110","000000000000000100","111111111111101010","000000000000001001","000000000000001001","000000000000001110","111111111111110110","000000000000000100","111111111111111011","000000000000000101","111111111111011010","000000000000000011","111111111111100001","111111111111101001","000000000000010001","000000000000001011","000000000000001010","111111111111100001","111111111111011000","000000000000010001","111111111111100100","000000000000000110","111111111111110111","000000000000000010","111111111110111100","111111111111111110","000000000000000111","111111111111111011","000000000000011111","111111111111110111","000000000000001000","000000000000001000","111111111111111110","111111111111111000","000000000000001000","111111111111111101","000000000000000100","000000000000010101","000000000000010101","111111111111100100","000000000000000001","111111111111100011","000000000000101001","111111111111011100","000000000000000011","000000000000010110","111111111111101101","000000000000000000","111111111111101101","000000000000011101","111111111111111101","111111111111101100","000000000000000010","111111111111110010","111111111111101101","111111111111110111","111111111111111111","000000000000011110","000000000000000000","000000000000001001","111111111111110100","000000000000011001","000000000000000101","111111111111111000","111111111111110000","111111111111111000","000000000000000010","000000000000010000","111111111111111110","111111111111111110","111111111111111000","111111111111111110","000000000000000011","000000000000001000","111111111111110101","111111111111101110","111111111111101111","111111111111111010","111111111111101101","000000000000110010","111111111111111101","000000000000000001","111111111111101011","000000000000001110"),
("000000000000001110","000000000000101100","000000000000111101","111111111111111110","000000000000000101","000000000000010111","000000000000000001","000000000000010010","111111111111000100","000000000000111111","111111111111011001","000000000000101101","111111111111010111","000000000000010111","111111111111111110","111111111111101110","111111111111111010","000000000000001101","111111111111110011","111111111111101000","000000000000001011","000000000000011100","000000000000001011","111111111111011101","000000000000001000","000000000000000100","000000000000011100","111111111111111001","111111111111010101","111111111111101110","000000000000010000","111111111111111111","000000000000000010","111111111111110011","111111111111110110","000000000000001000","000000000000001101","111111111111110101","000000000000001010","111111111111101010","000000000000001011","111111111111101001","111111111111001000","111111111111110010","000000000000000111","000000000000001000","111111111111001010","000000000000001100","000000000000011000","000000000000000000","111111111111100000","111111111111111101","000000000000010101","000000000000000011","111111111111110001","000000000000000011","111111111111011110","111111111111111111","000000000000011110","111111111111111011","111111111111110011","111111111111110101","111111111111110111","000000000000100001","111111111111110011","000000000000100100","111111111111110011","000000000000001010","111111111110010000","000000000000011110","000000000000001001","111111111111111010","000000000000100010","000000000000000010","000000000000000110","000000000000011011","000000000000010011","111111111111110110","111111111111110111","111111111111111010","000000000000010111","000000000000010111","000000000000001110","111111111111110111","111111111111110001","000000000000010110","000000000000101110","000000000000000111","000000000000001111","111111111111100011","111111111111111100","000000000000010010","000000000000001111","000000000000001000","000000000000001100","111111111111100101","000000000000101001","111111111111101011","111111111111001110","111111111111110001","000000000000011000","000000000000011110","000000000000000000","000000000000001111","111111111111011101","111111111111110100","000000000000001011","000000000000010000","111111111111110111","000000000000000111","000000000000000010","111111111111111110","000000000000000101","111111111111100000","111111111111011001","111111111111111011","111111111111011001","111111111111100101","000000000000000110","111111111111111010","111111111111111000","000000000000000000","111111111111100001","000000000000011001","111111111111110111","000000000000011111","111111111111100010","000000000000011111"),
("000000000000000000","000000000000100000","000000000000110100","000000000000001111","111111111111111110","000000000000011010","000000000000011101","111111111111101110","111111111111110110","000000000000111010","111111111111101011","000000000000010110","111111111111110111","000000000000001001","000000000000001011","111111111111010100","111111111111101011","111111111111101000","111111111111111100","111111111111101111","000000000000010000","000000000000011100","000000000000001111","111111111111011010","111111111111111000","111111111111111001","000000000000000110","111111111111101111","000000000000000000","111111111111111111","111111111111111111","000000000000001001","111111111111101111","000000000000000000","111111111111101011","000000000000010100","111111111111110000","000000000000000000","000000000000010010","111111111111110110","111111111111111001","111111111111110101","111111111111011000","000000000000000001","111111111111111011","111111111111110111","111111111111010111","000000000000000000","111111111111111111","111111111111110001","000000000000000110","000000000000010000","000000000000000101","111111111111110011","111111111111110100","000000000000000001","000000000000001100","000000000000000011","000000000000000011","111111111111111111","111111111111110111","000000000000010011","111111111111100101","000000000000010101","111111111111111000","000000000000010001","111111111111110010","000000000000000101","111111111110011110","000000000000010100","111111111111110001","111111111111101011","111111111111111110","000000000000000100","111111111111101100","000000000000010001","111111111111111001","000000000000000110","000000000000000011","111111111111111111","000000000000010000","111111111111111010","000000000000001110","111111111111100011","111111111111111010","000000000000001000","000000000000100111","000000000000001100","000000000000010111","111111111111110010","000000000000001000","000000000000010101","111111111111111011","000000000000001111","000000000000010010","111111111111111000","000000000000000000","111111111111101110","111111111111001111","111111111111101100","000000000000001110","000000000000100001","000000000000001100","000000000000001111","111111111111100000","111111111111111110","000000000000001101","000000000000000001","111111111111111100","000000000000001000","000000000000000010","111111111111011100","000000000000011011","000000000000000000","111111111111111110","000000000000010010","111111111111111110","111111111111110110","000000000000010011","111111111111011011","111111111111100001","111111111111101011","000000000000000000","000000000000011111","111111111111111110","111111111111110000","111111111111100000","000000000000000010"),
("000000000000000100","000000000000000000","000000000000101100","000000000000000011","000000000000001110","000000000000011011","111111111111110100","111111111111100001","111111111111101010","000000000001000000","111111111111100000","000000000000010101","111111111111100100","111111111111110010","000000000000010001","000000000000000000","000000000000001000","000000000000001000","000000000000000000","111111111111100010","111111111111111010","000000000000100111","000000000000001100","111111111111110110","111111111111111110","111111111111100100","000000000000100111","111111111111110110","111111111111110010","000000000000001010","111111111111110100","111111111111011111","111111111111110010","111111111111101011","111111111111111010","000000000000010100","111111111111111101","111111111111101111","111111111111111111","000000000000001010","111111111111110100","000000000000010010","111111111111010000","000000000000000000","111111111111111110","000000000000010011","111111111111101000","000000000000000001","000000000000100001","111111111111110111","000000000000010000","111111111111111111","000000000000000110","111111111111111010","000000000000000011","111111111111101111","111111111111111010","111111111111101111","000000000000010001","111111111111111111","111111111111101100","000000000000001010","111111111111111111","000000000000000101","000000000000000000","000000000000100100","000000000000000001","000000000000000011","111111111110011110","000000000000101010","111111111111110000","111111111111111001","000000000000000000","000000000000000000","111111111111110010","000000000000010100","000000000000001000","000000000000000010","111111111111110111","111111111111110100","000000000000011111","111111111111111001","000000000000001100","111111111111000011","000000000000001111","000000000000001000","000000000000001010","000000000000100100","000000000000100001","000000000000100010","000000000000000010","000000000000000100","000000000000010101","000000000000001010","000000000000011010","000000000000000000","000000000000000000","111111111111110110","111111111111111000","111111111111111100","000000000000100011","000000000000101010","000000000000011000","000000000000000000","111111111111101011","000000000000001101","000000000000000001","111111111111101101","111111111111110000","111111111111111100","111111111111111010","111111111111011110","000000000000011001","111111111111111110","000000000000000011","000000000000000000","111111111111110001","111111111111111001","000000000000000101","111111111111101100","111111111111010010","111111111111110001","111111111111111010","000000000000110000","111111111111111111","000000000000100000","111111111111111110","000000000000011001"),
("000000000000000111","111111111111100010","000000000000010010","111111111111101110","111111111111110100","000000000000001001","000000000000001000","111111111111110001","111111111111101011","000000000000101111","111111111110101001","000000000000011100","111111111111011110","111111111111100010","000000000000001110","111111111111110011","000000000000100001","111111111111011110","111111111111011110","000000000000000100","111111111111101011","000000000000000111","111111111111100111","000000000000000111","000000000000010011","111111111111011011","000000000000010011","111111111111101101","000000000000001001","000000000000001110","111111111111110000","111111111111011101","000000000000000111","000000000000000110","111111111111110010","111111111111110101","000000000000010001","111111111111110110","000000000000010001","000000000000000000","000000000000000101","000000000000000101","111111111111011110","000000000000000110","000000000000100011","000000000000101101","111111111111001100","111111111111110110","000000000000010011","111111111111111010","000000000000011101","000000000000010101","000000000000010110","111111111111100000","111111111111111110","000000000000001001","000000000000100000","000000000000000000","000000000000001110","111111111111111100","000000000000000001","000000000000100011","000000000000011010","000000000000000000","000000000000001110","000000000000001101","000000000000000101","000000000000010111","111111111111010010","000000000000010100","111111111111101001","111111111111100100","000000000000000100","111111111111110100","000000000000000000","000000000000001101","000000000000000111","111111111111100111","000000000000000100","111111111111110111","000000000000010011","000000000000011111","000000000000001010","111111111110111000","111111111111100001","000000000000010010","000000000000011011","000000000000001111","000000000000100001","000000000000010011","000000000000101010","111111111111101010","000000000000011100","111111111111110010","111111111111111101","000000000000001100","000000000000001111","111111111111111100","000000000000100010","111111111111110010","000000000000010001","000000000000101111","000000000000001000","111111111111111010","111111111111100100","111111111111110110","000000000000001101","000000000000001110","000000000000001011","000000000000011000","111111111111110001","111111111111101000","000000000000010001","111111111111101111","111111111111101001","000000000000001110","000000000000001100","111111111111101000","000000000000001000","111111111111101110","111111111111111011","111111111111110100","111111111111101000","000000000000101010","000000000000101111","000000000000100111","111111111111101001","000000000000010100"),
("000000000000010111","111111111110111000","000000000000000111","111111111111100110","111111111111110010","111111111111110000","111111111111101111","111111111111111101","111111111111110100","000000000000100111","111111111110011011","000000000000100000","111111111111011001","111111111111100100","000000000000011011","111111111111110110","000000000000011101","111111111111101101","111111111111101000","000000000000000111","111111111111100000","111111111111110001","111111111111100101","111111111111111101","000000000000000010","111111111111101111","000000000000011110","111111111111010000","111111111111110100","000000000000010101","000000000000000010","111111111111100111","000000000000001111","000000000000000001","111111111111111111","000000000000001101","000000000000001101","111111111111111000","000000000000100100","111111111111111101","111111111111110100","000000000000001011","111111111111100000","000000000000001000","000000000000011011","000000000000010111","111111111111011010","000000000000010000","000000000000001101","111111111111110001","000000000000101101","000000000000110000","000000000000001110","111111111111110010","111111111111100111","111111111111111010","111111111111111110","111111111111110111","111111111111111011","111111111111101100","111111111111100111","000000000000011000","000000000000101011","111111111111111011","000000000000010110","000000000000100000","000000000000010010","000000000000010001","111111111111100000","000000000000011010","111111111111110000","111111111111010000","000000000000000110","000000000000000111","000000000000000100","000000000000100010","000000000000000000","111111111111011101","000000000000001111","000000000000000010","000000000000001100","000000000000100000","111111111111101101","111111111111011001","111111111111110001","000000000000100100","000000000000100000","000000000000100001","000000000000010010","000000000000010110","000000000000010111","000000000000010010","000000000000000001","000000000000001001","000000000000001000","111111111111110111","000000000000011110","000000000000011111","000000000000010000","111111111111110001","111111111111111101","000000000000011001","111111111111101101","111111111111110100","000000000000000001","000000000000010100","111111111111110000","111111111111101010","000000000000001000","000000000000101111","000000000000000010","111111111111011111","000000000000001100","000000000000100100","000000000000001001","111111111111111101","111111111111110010","111111111111101001","000000000000001100","111111111111011011","111111111111010101","111111111111111001","111111111111110110","000000000000000000","000000000000100101","000000000000001110","111111111111101000","000000000000001000"),
("000000000000100010","111111111110101001","111111111111110110","111111111111111000","111111111111110101","000000000000001110","111111111111110001","000000000000001101","000000000000000000","111111111111100111","111111111110101000","000000000000100100","111111111111000101","111111111111110100","111111111111011111","000000000000010111","000000000000011001","111111111111111010","111111111111000011","000000000000000110","111111111111100101","111111111111111111","111111111111011111","000000000000001110","000000000000100111","000000000000010111","000000000000100011","111111111111011010","000000000000010010","000000000000001111","111111111111110011","111111111111110100","000000000000010111","111111111111111110","111111111111100101","000000000000011110","111111111111101110","000000000000011100","000000000000011111","111111111111111000","111111111111101011","111111111111111100","111111111111101010","111111111111110101","000000000000010100","111111111111110001","000000000000000101","000000000000111010","000000000000010111","000000000000001001","000000000000100000","000000000000010110","111111111111111000","111111111111100101","111111111111111110","111111111111101100","000000000000000101","111111111111011010","000000000000000001","111111111111111000","111111111111110011","000000000000010101","000000000000011110","000000000000001011","000000000000100001","000000000000001000","000000000000000000","111111111111111111","111111111111100111","111111111111111110","000000000000010111","111111111111010101","000000000000001100","111111111111110001","000000000000010011","000000000000100101","000000000000010001","000000000000000001","111111111111101101","000000000000010100","000000000000010111","000000000000011011","111111111111101001","111111111111010000","111111111111110011","000000000000011001","000000000000101001","000000000000000111","000000000000000100","000000000000011110","000000000000010110","000000000000001110","111111111111101101","000000000000000000","111111111111110111","000000000000001011","000000000000001000","000000000000000001","000000000000101001","111111111111100001","111111111111111101","000000000000011000","000000000000001110","000000000000001100","111111111111110110","000000000000011111","000000000000000000","111111111111100001","000000000000001001","000000000000010011","111111111111111001","111111111111011001","000000000000011101","000000000000010001","000000000000000000","000000000000000000","111111111111110101","111111111111111001","000000000000101010","000000000000000101","111111111111110000","000000000000100010","111111111111100011","111111111111001011","000000000000100101","000000000000010011","111111111111101010","000000000000000000"),
("000000000000100100","111111111111000101","111111111111101101","000000000000010000","111111111111111011","000000000000001011","111111111111110010","111111111111110101","000000000000100000","111111111111001000","111111111111100110","000000000000000011","111111111111001111","000000000000001011","111111111111101001","000000000000010000","000000000000001101","000000000000010001","111111111111011101","111111111111111010","111111111111101110","111111111111111111","111111111111001010","000000000000001101","111111111111110111","000000000000101110","000000000000001111","111111111111111000","000000000000010101","000000000000011100","000000000000000100","111111111111111010","000000000000011100","111111111111111010","111111111111101100","000000000000010111","000000000000001000","000000000000001110","000000000000100011","111111111111111100","111111111111011011","000000000000000100","000000000000011001","111111111111111101","000000000000110011","111111111111111001","000000000000011000","000000000000101101","000000000000010101","000000000000001111","111111111111111111","000000000000010000","111111111111101001","000000000000001101","111111111111111101","111111111111111000","000000000000010000","111111111111100111","111111111111101101","000000000000001001","000000000000010111","000000000000100000","111111111111110111","000000000000010101","000000000000101000","000000000000000111","111111111111110100","000000000000011110","000000000000001011","111111111111001010","000000000000100101","111111111111111000","000000000000001100","111111111111111100","000000000000101011","000000000000010100","111111111111111100","000000000000010111","111111111111100101","111111111111111101","000000000000010110","000000000000100101","111111111111101010","000000000000000111","000000000000011001","000000000000000011","000000000000001000","000000000000011011","111111111111101100","000000000000100010","111111111111110001","000000000000001001","111111111111110010","111111111111101100","111111111111111000","000000000000101101","000000000000011100","000000000000000000","000000000000110011","111111111111111000","111111111111110100","000000000000000111","000000000000010110","000000000000010000","000000000000010011","000000000000011010","000000000000000101","111111111111101100","000000000000100010","111111111111100101","000000000000000011","111111111111001111","000000000000011000","000000000000011011","000000000000000101","111111111111101110","000000000000010111","111111111111101010","000000000000101010","111111111111111001","111111111111110100","000000000000010111","111111111111101100","111111111110011000","000000000000001010","111111111111101110","111111111111110100","000000000000011011"),
("000000000000101110","111111111111100101","111111111111110001","111111111111111000","111111111111110010","000000000000001011","111111111111101100","111111111111110101","000000000000010100","111111111111101110","111111111111111111","111111111111110110","000000000000001001","000000000000110110","111111111111111010","111111111111101001","000000000000000000","000000000000000000","111111111111110110","111111111111101010","000000000000001001","000000000000010001","111111111111010001","000000000000001111","111111111111110101","000000000000001100","111111111111100101","111111111111111111","000000000000100011","000000000000000110","000000000000010100","000000000000010010","000000000000010010","111111111111111100","000000000000010101","000000000000110101","000000000000000101","000000000000000111","111111111111111100","000000000000000010","111111111111110100","000000000000011110","000000000000101011","000000000000001001","000000000000001011","111111111111101110","000000000000111010","000000000000000110","111111111111111110","000000000000001111","000000000000000110","000000000000000101","111111111111110101","000000000000000001","000000000000011110","111111111111111100","000000000000011001","111111111111101010","111111111111111010","000000000000000000","000000000000001111","000000000000010101","111111111111111101","000000000000000001","000000000001001001","111111111111111110","000000000000011001","000000000000000011","000000000000001101","111111111111011101","000000000000011011","111111111111111011","111111111111111010","000000000000011000","000000000000110100","000000000000001100","000000000000000100","000000000000011001","111111111111100100","111111111111110000","111111111111111010","000000000000000010","111111111111011001","000000000000110010","111111111111111010","111111111111101101","000000000000000000","000000000000010010","111111111111101010","000000000000011111","111111111111100111","000000000000010000","000000000000000001","000000000000000111","111111111111100110","000000000000100101","000000000000000111","000000000000010110","000000000000001011","111111111111111001","000000000000000001","111111111111110000","000000000000011011","000000000000100110","111111111111111111","111111111111110101","000000000000001100","111111111111100111","000000000000001011","111111111111110110","000000000000011011","111111111111110100","000000000000100100","000000000000000101","111111111111101111","111111111111111001","000000000000000000","111111111111101101","000000000000011101","111111111111111011","111111111111110111","111111111111111001","000000000000011010","111111111110110010","000000000000001011","111111111111101000","111111111111101010","000000000000001111"),
("000000000000001100","000000000000000001","000000000000001111","111111111111110101","000000000000000110","000000000000011110","000000000000000111","000000000000010011","000000000000011100","111111111111101101","111111111111011011","111111111111110111","111111111111111111","000000000000011010","000000000000000010","111111111111100111","111111111111011111","000000000000010110","111111111111101111","111111111111010101","111111111111101100","000000000000001000","111111111111000111","000000000000010110","111111111111101111","000000000000001010","111111111111111001","000000000000000011","000000000000010011","111111111111011111","000000000000000111","000000000000001010","111111111111100000","000000000000010001","000000000000000110","000000000000110001","000000000000000001","000000000000011110","000000000000000111","111111111111110100","111111111111111001","000000000000100111","000000000000110001","000000000000000001","000000000000011000","111111111111101101","000000000000001001","000000000000100101","111111111111110110","000000000000001011","000000000000010101","000000000000001110","111111111111110101","000000000000000110","000000000000011001","000000000000011000","000000000000001101","000000000000000010","111111111111111010","111111111111101101","000000000000001010","000000000000001111","111111111111110001","000000000000010100","000000000000111000","000000000000000000","111111111111110111","000000000000011001","111111111111110010","111111111111011100","000000000000100101","111111111111111111","111111111111010111","111111111111111101","000000000000100110","111111111111111111","111111111111111011","111111111111111001","000000000000001000","111111111111101101","000000000000010001","000000000000000010","111111111111101011","000000000000101011","000000000000000001","111111111111111101","111111111111110101","111111111111110101","000000000000000001","111111111111101101","000000000000001100","111111111111111101","111111111111111110","000000000000000000","000000000000000100","000000000000010101","111111111111100011","000000000000101101","000000000000000000","000000000000001111","111111111111101100","111111111111110111","111111111111110101","000000000000010011","000000000000000011","000000000000000001","000000000000001100","000000000000001100","000000000000000100","111111111111110110","000000000000001110","111111111111010010","000000000000001110","000000000000100100","000000000000000011","000000000000000110","000000000000000110","111111111111001111","000000000000001111","111111111111111011","111111111111101100","111111111111110110","000000000000011100","111111111111100011","000000000000001111","111111111111110110","111111111111111000","000000000000010111"),
("000000000000100101","111111111111110000","000000000000001000","111111111111111110","000000000000100101","000000000000001011","000000000000001000","000000000000010000","000000000000100011","111111111111110001","111111111111010110","111111111111011101","111111111111110010","000000000000010001","000000000000000001","111111111111110000","000000000000001000","111111111111111000","000000000000000110","111111111111101111","111111111111101110","000000000000010001","111111111111111001","000000000000001100","111111111111101011","000000000000010000","111111111111111101","000000000000001001","111111111111110101","111111111111101010","000000000000000111","000000000000100101","111111111111100111","000000000000001000","000000000000001111","000000000000101100","111111111111100110","000000000000000011","000000000000010100","000000000000001100","111111111111111000","111111111111101101","000000000000011101","000000000000100000","000000000000010100","000000000000001110","000000000000001101","000000000000000100","000000000000001101","111111111111111100","000000000000100000","111111111111011100","000000000000001100","000000000000000011","000000000000001111","000000000000000000","000000000000011101","111111111111101010","000000000000000111","000000000000001110","111111111111111100","000000000000001001","111111111111111000","000000000000000010","000000000000011000","111111111111110101","000000000000001101","111111111111110100","111111111111101111","111111111111110011","000000000000000000","111111111111111001","111111111111011010","000000000000000111","000000000000010100","000000000000001100","000000000000010010","111111111111111101","000000000000100000","000000000000010000","000000000000001010","000000000000000000","111111111111111110","000000000000001001","111111111111111101","000000000000101010","111111111111100011","111111111111111001","000000000000011100","111111111111111110","000000000000000011","000000000000001000","111111111111100000","111111111111011110","111111111111111000","000000000000010111","111111111111011111","000000000000101111","111111111111111010","000000000000110000","000000000000000010","111111111111100111","111111111111110011","000000000000000001","111111111111111101","000000000000000111","000000000000010010","000000000000100110","000000000000011100","000000000000000111","000000000000001011","111111111111100100","000000000000000010","000000000000001111","000000000000000000","111111111111110001","000000000000000101","111111111111110101","111111111111111100","000000000000001001","111111111111111010","111111111111101010","000000000000110111","000000000000000110","111111111111111001","000000000000000101","111111111111011111","000000000000011111"),
("000000000000001001","000000000000001100","000000000000000011","111111111111110010","000000000000001001","111111111111110111","111111111111111111","111111111111110010","000000000000001011","111111111111110011","000000000000000010","000000000000000000","111111111111111111","000000000000001001","000000000000001010","111111111111011100","111111111111111000","111111111111110011","111111111111101111","111111111111111011","000000000000000000","000000000000010011","111111111111101111","111111111111111101","111111111111101101","000000000000001000","111111111111111111","000000000000000000","111111111111111111","111111111111110000","111111111111111010","000000000000010101","000000000000001010","111111111111111001","111111111111100111","000000000000011010","111111111111110101","000000000000001111","111111111111111001","000000000000011000","000000000000010000","111111111111100001","000000000000001010","000000000000100000","000000000000011000","000000000000001110","111111111111111100","000000000000010110","000000000000000001","000000000000001100","000000000000000110","111111111111100100","111111111111111110","000000000000001001","000000000000011100","000000000000001010","000000000000001111","111111111111110010","000000000000010111","111111111111110011","111111111111110100","111111111111101111","111111111111111000","000000000000000100","000000000000110001","000000000000000111","000000000000000000","111111111111110101","111111111111111010","111111111111110100","000000000000001100","111111111111110010","111111111111110011","000000000000001000","000000000000011110","111111111111111001","000000000000000111","000000000000000111","000000000000001100","000000000000000001","111111111111110011","111111111111111110","000000000000001100","000000000000001111","111111111111111010","000000000000100110","000000000000000101","111111111111111010","000000000000001110","111111111111100011","000000000000001110","000000000000000000","111111111111011101","111111111111010100","000000000000000010","000000000000010001","111111111111101111","000000000000011111","000000000000000001","000000000000010010","111111111111110110","111111111111111111","111111111111110110","000000000000000111","111111111111110100","000000000000000011","000000000000010001","111111111111111100","000000000000100110","111111111111111110","000000000000011000","111111111111101000","000000000000000110","000000000000000110","000000000000011001","111111111111011111","111111111111111100","000000000000001011","000000000000000011","000000000000001010","111111111111110010","000000000000000001","000000000000011010","000000000000010100","000000000000000111","000000000000000110","111111111111010101","000000000000000101"),
("111111111111110011","000000000000000001","111111111111101111","000000000000001010","111111111111011111","111111111111111111","000000000000001101","111111111111110010","000000000000000111","111111111111110000","000000000000000011","000000000000000101","111111111111111000","000000000000011110","000000000000000000","111111111111111001","000000000000000101","111111111111110011","111111111111010111","000000000000000000","111111111111101000","000000000000001101","111111111111111100","111111111111111001","111111111111011110","111111111111101000","000000000000001010","000000000000000011","111111111111101101","111111111111011010","000000000000000101","000000000000011001","000000000000000101","000000000000011001","111111111111101101","000000000000001111","000000000000000100","111111111111111000","000000000000000010","000000000000000100","111111111111101000","000000000000000101","000000000000011100","000000000000101011","000000000000011100","000000000000001100","000000000000010101","111111111111111111","000000000000000011","111111111111111110","000000000000001100","000000000000010000","000000000000000101","111111111111101111","000000000000010000","000000000000011101","000000000000000111","000000000000011001","000000000000011111","111111111111111010","000000000000000000","111111111111110100","000000000000010000","000000000000010001","111111111111101110","000000000000000000","111111111111011010","111111111111110110","111111111111111010","111111111111111001","111111111111111100","111111111111110100","111111111111111000","000000000000100001","111111111111111110","111111111111111100","000000000000010000","000000000000001000","000000000000001011","000000000000000110","111111111111111010","000000000000011010","111111111111111010","000000000000000100","111111111111111000","000000000000111000","000000000000011101","000000000000010100","000000000000100000","111111111111100001","000000000000000010","111111111111110001","111111111111011100","111111111111101101","000000000000000110","111111111111111111","111111111111111011","000000000000011000","000000000000011110","000000000000100110","111111111111110000","000000000000000000","000000000000000110","000000000000001001","111111111111101111","000000000000000110","000000000000100000","000000000000011001","000000000000001111","000000000000001011","000000000000001110","111111111111101000","000000000000001011","000000000000000110","000000000000011001","111111111111101110","000000000000001101","000000000000010001","111111111111111011","111111111111111000","000000000000001001","111111111111111101","111111111111110101","111111111111111101","000000000000010000","111111111111111011","111111111111100100","000000000000011001"),
("111111111111111101","111111111111111011","111111111111100010","000000000000001111","111111111111100010","111111111111110011","000000000000010100","111111111111110000","111111111111110000","111111111111110111","111111111111110101","111111111111101010","000000000000001000","000000000000000101","111111111111111011","111111111111111000","111111111111111100","000000000000000001","111111111111101111","111111111111101001","111111111111010111","111111111111110100","111111111111001101","000000000000000011","000000000000000100","000000000000010011","000000000000010010","000000000000000000","111111111111111001","111111111111100111","111111111111111000","000000000000001101","000000000000100011","000000000000101100","111111111111101110","111111111111011011","111111111111101011","111111111111101000","111111111111110011","111111111111111010","111111111111111001","000000000000100110","111111111111111011","000000000000100111","000000000000010001","111111111111110100","000000000000010011","000000000000011011","111111111111111100","000000000000000011","111111111111111011","000000000000010011","111111111111110011","111111111111111010","111111111111110011","000000000000001110","000000000000001001","111111111111111010","000000000000010111","000000000000001001","111111111111110110","111111111111110100","111111111111110101","000000000000001101","111111111111010011","000000000000001101","111111111111010111","111111111111110001","111111111111110000","111111111111101011","111111111111111101","111111111111011010","111111111111101000","111111111111111101","111111111111111000","111111111111111011","000000000000010000","000000000000010111","111111111111110101","111111111111111010","111111111111101110","000000000000010101","111111111111110100","000000000000000110","000000000000001001","000000000000100000","000000000000010011","000000000000001001","000000000000011010","000000000000000001","111111111111101010","111111111111100101","000000000000000010","111111111111101101","000000000000010110","000000000000001001","111111111111101000","000000000000101010","000000000000000101","000000000000001101","111111111111111011","000000000000010010","000000000000001100","111111111111110110","111111111111011110","000000000000001001","000000000000011000","000000000000101111","000000000000011111","000000000000100110","000000000000010001","000000000000010111","000000000000010111","000000000000010101","000000000000010001","000000000000011100","000000000000000001","000000000000010010","000000000000010011","000000000000000100","000000000000000001","000000000000000000","111111111111011101","111111111111101101","000000000000011101","000000000000000010","111111111111011010","000000000000001110"),
("111111111111100101","111111111111111100","000000000000001001","111111111111111100","000000000000000000","111111111111111110","000000000000100101","111111111111110010","111111111111111101","111111111111111010","000000000000001001","111111111111101000","111111111111111100","111111111111111001","000000000000100010","111111111111101000","000000000000001000","000000000000000101","111111111111101010","111111111111100001","111111111111110101","000000000000000011","111111111111010000","000000000000000000","000000000000000010","111111111111110110","000000000000000111","111111111111111110","111111111111111100","111111111111010101","000000000000000100","000000000000000111","111111111111111100","000000000000001101","111111111111101111","111111111111011111","111111111111110001","000000000000000111","000000000000000111","000000000000000101","000000000000000101","000000000000100101","000000000000000000","111111111111110110","000000000000010111","000000000000000010","000000000000100100","000000000000000000","000000000000011000","000000000000000000","111111111111110100","000000000000010100","111111111111111100","000000000000000101","111111111111110111","000000000000100100","111111111111111010","111111111111101001","000000000000011001","111111111111110100","111111111111110111","000000000000000001","000000000000010000","000000000000001001","111111111111000110","000000000000000001","111111111111101100","111111111111110101","111111111111110101","111111111111100100","111111111111110111","111111111111100011","111111111111011110","111111111111010110","000000000000010101","111111111111111111","111111111111111111","000000000000100011","000000000000011011","000000000000001011","000000000000000000","000000000000010110","111111111111110110","000000000000010000","111111111111110111","000000000000011001","000000000000100011","000000000000001000","000000000000010100","000000000000010010","111111111111101011","111111111111101000","111111111111111000","000000000000001001","111111111111111101","000000000000000000","111111111111100111","000000000000001101","000000000000000110","000000000000101110","111111111111101111","000000000000010111","111111111111110101","111111111111111101","111111111111100111","000000000000001010","000000000000000000","000000000000100011","000000000000010011","000000000000000110","000000000000011000","000000000000011101","111111111111111111","111111111111110101","000000000000001011","000000000000000110","111111111111110000","000000000000001001","000000000000010011","000000000000000010","000000000000000100","111111111111111111","111111111111001111","111111111111111111","000000000000001010","111111111111101110","111111111111010000","111111111111111000"),
("111111111111000010","000000000000100011","000000000000001001","111111111111111101","000000000000010101","111111111111110110","000000000000010111","111111111111101001","000000000000000000","000000000000000011","000000000000000100","000000000000000000","111111111111110001","111111111111010111","000000000000101011","000000000000001000","000000000000010111","111111111111100000","000000000000000001","111111111111100100","000000000000000110","000000000000010111","111111111111100111","000000000000100010","000000000000000101","111111111111110101","000000000000011011","000000000000000101","111111111111101100","111111111111001101","111111111111100101","000000000000010000","000000000000000000","111111111111100001","000000000000001101","111111111111010011","111111111111111111","000000000000000001","111111111111101010","111111111111100101","111111111111111000","000000000000100110","000000000000000110","111111111111110010","000000000000000010","111111111111111101","000000000000000011","111111111111111110","000000000000000011","000000000000000111","000000000000010000","111111111111101010","111111111111110101","111111111111111100","111111111111101010","111111111111110111","111111111111100011","111111111111111111","000000000000000011","000000000000001110","111111111111110000","111111111111111100","000000000000001011","000000000000100001","111111111111000101","000000000000010100","111111111111000110","111111111111101010","111111111111110001","111111111111110110","000000000000010100","111111111111101110","111111111111100000","111111111111111011","000000000000010000","111111111111110010","000000000000000001","000000000000001001","000000000000100010","111111111111111001","000000000000001100","000000000000001100","111111111111111111","000000000000011101","111111111111110111","000000000000001001","000000000000110100","000000000000001011","111111111111110110","000000000000010010","111111111111111101","111111111111111110","111111111111110111","000000000000010110","000000000000000000","111111111111110100","000000000000001100","000000000000001000","111111111111111001","000000000000010111","000000000000010111","000000000000101001","000000000000001001","111111111111011010","000000000000000000","000000000000010100","000000000000000010","000000000000101101","000000000000001110","000000000000010100","000000000000010101","000000000000011111","111111111111111111","111111111111101010","000000000000010111","000000000000001111","000000000000001011","111111111111101001","111111111111110100","000000000000000101","111111111111100000","111111111111110011","000000000000001001","000000000000000011","000000000000010001","000000000000000110","111111111111011000","000000000000000000"),
("111111111110111010","000000000000010011","111111111111111111","111111111111111100","000000000000011000","000000000000000001","000000000000010011","000000000000001001","111111111111111101","111111111111111111","111111111111101111","000000000000000111","111111111111011100","111111111110111111","000000000000001111","111111111111110100","000000000000001001","111111111111011110","111111111111011110","111111111111111010","000000000000001000","000000000000100110","000000000000001001","000000000000101011","000000000000010101","111111111111101101","111111111111111111","111111111111111000","111111111111101111","111111111111001001","111111111111011010","111111111111111101","111111111111111101","111111111111110001","111111111111111011","111111111111110100","111111111111101100","111111111111100011","111111111111110001","111111111111100011","111111111111111001","111111111111101101","000000000000100110","111111111111110110","000000000000000011","111111111111111110","111111111111111001","000000000000000111","111111111111101010","111111111111111111","000000000000011000","000000000000000010","000000000000001101","000000000000010001","111111111111100010","000000000000010001","111111111111010100","000000000000000011","000000000000000110","000000000000000111","000000000000001110","000000000000001001","111111111111011110","000000000000010000","111111111110111111","000000000000010111","111111111111001010","111111111111110111","111111111111011010","111111111111101111","000000000000001011","111111111111100100","111111111111001010","111111111111011110","111111111111111100","111111111111111101","000000000000000110","000000000000001000","000000000000000101","000000000000010101","000000000000001010","111111111111111110","000000000000010010","000000000000001100","111111111111111100","111111111111100110","000000000000011111","111111111111101101","000000000000000011","000000000000010000","111111111111110101","111111111111110111","111111111111111111","000000000000001111","000000000000010011","111111111111100110","000000000000001110","000000000000011011","111111111111010100","111111111111101101","000000000000000011","000000000000100010","000000000000010001","111111111111100100","000000000000010100","000000000000001111","000000000000001101","000000000000010101","000000000000010101","111111111111111111","111111111111101111","000000000000100001","000000000000010000","111111111111010101","111111111111101111","000000000000001011","111111111111111010","111111111111011110","111111111111101110","111111111111110110","111111111111011010","000000000000100001","111111111111111010","111111111111111001","111111111111110111","000000000000000111","111111111111010101","111111111111101001"),
("111111111110111011","000000000000100111","111111111111100111","111111111111100001","000000000000000001","000000000000010010","000000000000100010","000000000000000101","111111111111110111","000000000000000001","111111111111101001","111111111111111001","111111111111111111","111111111111010101","111111111111111111","111111111111111110","000000000000000110","111111111111110011","111111111111010101","111111111111110001","000000000000000011","000000000000010000","000000000000000000","000000000000100100","111111111111111111","000000000000010110","111111111111100101","111111111111101111","000000000000100011","000000000000000100","111111111111100111","000000000000010110","000000000000001100","111111111111110111","000000000000001000","111111111111111011","111111111111011011","111111111111011010","111111111111100011","111111111111010110","111111111111110111","111111111111111010","000000000000011111","111111111111101101","111111111111111000","000000000000001001","000000000000100100","000000000000011100","111111111111011111","000000000000000010","000000000000011101","111111111111110010","000000000000011010","000000000000001111","111111111111101101","111111111111100101","111111111111011101","111111111111011101","111111111111111010","111111111111111011","111111111111101001","111111111111011011","111111111111001111","111111111111111010","111111111111010100","000000000000000111","111111111111001011","000000000000110010","111111111111110011","111111111111110000","000000000000011110","111111111111000111","111111111111101000","111111111111100100","000000000000000111","000000000000000101","111111111111101001","111111111111010001","111111111111111010","000000000000100101","000000000000000011","000000000000001110","000000000000011100","000000000000000100","111111111111110011","111111111111101110","000000000000100101","000000000000001000","000000000000000010","000000000000100001","111111111111101011","111111111111110110","000000000000011010","000000000000011111","111111111111100000","111111111110111110","000000000000001011","000000000000001111","111111111110101110","111111111111000100","000000000000101011","000000000000101000","000000000000011011","111111111111011000","000000000000100010","000000000000100100","111111111111101110","000000000000010001","111111111111111001","111111111111110111","111111111111010111","000000000000010000","000000000000011110","111111111111100100","111111111111010110","000000000000101011","000000000000100011","111111111111011001","111111111111101100","111111111111101111","111111111111001101","000000000000000011","111111111111110000","111111111111110010","000000000000101011","000000000000010100","111111111111111011","111111111111100001"),
("111111111110110011","000000000000000000","111111111111111101","111111111111101110","111111111111011111","000000000000001110","000000000000010000","111111111111110111","000000000000011001","000000000000101001","000000000000000111","000000000000011110","111111111111011011","111111111111100001","111111111111101010","000000000000001000","000000000000011101","111111111111111001","111111111111110000","000000000000000001","000000000000001011","111111111111101010","000000000000010000","000000000000001100","000000000000001000","000000000000011110","111111111111101001","111111111111101100","111111111111111111","111111111111111001","111111111111101001","000000000000001000","000000000000001000","111111111111101011","111111111111111001","111111111111101001","111111111111011011","111111111111111101","111111111111101010","111111111111000000","000000000000010001","111111111111101000","000000000000000100","111111111111110100","111111111111101100","111111111111110100","000000000000011000","000000000000100000","111111111111011001","111111111111001101","000000000000010110","111111111111110001","000000000000010101","111111111111111111","000000000000000101","000000000000001010","111111111111011001","111111111111100010","000000000000000000","000000000000001101","111111111111100001","111111111111101111","111111111111101100","111111111111100010","111111111111110010","111111111111110110","111111111111000011","000000000000001000","000000000001000101","000000000000000011","000000000000000111","111111111111010000","111111111110111110","000000000000010110","111111111111111001","000000000000100110","111111111111110111","111111111111111000","111111111111111110","000000000000011000","111111111111011011","111111111111010000","000000000000001010","111111111111101111","111111111111101011","111111111111100111","000000000000001101","111111111111100011","111111111111100011","111111111111110111","111111111111110000","111111111111011010","000000000000101010","000000000000011100","111111111111010010","111111111110111111","000000000000110101","000000000000010101","111111111110101111","111111111111011110","000000000000001001","111111111111111010","111111111111001011","111111111111011000","000000000000100111","000000000000011111","111111111111100010","000000000000001110","111111111111110000","111111111111110101","111111111111001111","111111111111111111","111111111111111001","111111111111101010","111111111111100101","000000000000011110","000000000000101100","111111111111110110","000000000000000011","111111111111111111","111111111110110101","000000000000010011","000000000000100011","111111111111110001","000000000000011110","000000000000000110","000000000000000001","111111111111011101"),
("111111111110111010","000000000000001011","000000000000010000","111111111111111010","111111111111111110","000000000000000010","000000000000000111","000000000000100111","000000000000010010","000000000000100011","111111111111110100","000000000000001001","111111111111011110","000000000000010101","111111111111011111","000000000000011001","000000000000001111","000000000000001011","111111111111101101","000000000000011100","000000000000001011","111111111111101110","111111111111111100","111111111111111000","111111111111101111","111111111111110100","000000000000000010","111111111111111001","000000000000001101","000000000000000000","111111111111111111","111111111111100110","111111111111101001","111111111111100011","000000000000011100","111111111111011111","000000000000001010","000000000000010110","111111111111100010","111111111111010011","111111111111010101","111111111111101110","000000000000001011","111111111111100100","111111111111100010","111111111111100111","000000000000000111","000000000000001000","111111111111111010","111111111111001101","111111111111111111","000000000000001000","111111111111110001","111111111111110110","000000000000001011","000000000000100011","111111111111011011","111111111111111000","111111111111011010","000000000000010100","111111111111011010","000000000000000011","000000000000010101","111111111111011011","111111111111100110","111111111111011100","111111111111110100","111111111111111010","000000000000101100","111111111111101101","111111111111101111","111111111111111011","111111111111101100","000000000000001100","111111111111011110","111111111111111110","000000000000000110","111111111111010111","000000000000001010","000000000000011111","111111111111100111","111111111111101100","000000000000100001","000000000000001110","111111111111101101","111111111111111111","000000000000000001","111111111111011111","111111111111000011","111111111111110001","111111111111001010","111111111111110001","111111111111110110","000000000000000001","111111111111111100","111111111111101011","000000000000101010","000000000000010111","111111111111010110","111111111111101010","000000000000011100","111111111111101101","111111111111001111","111111111111110100","000000000000010110","000000000000001010","000000000000001001","111111111111111001","000000000000000000","111111111111110111","111111111111110110","111111111111100101","111111111111011011","111111111111110100","000000000000010000","111111111111110111","111111111111101011","000000000000000001","111111111111110100","111111111111001111","111111111111011000","000000000000100110","000000000000001111","111111111111100011","000000000000011111","111111111111111000","000000000000000000","111111111111110111"),
("111111111111100101","111111111111001011","111111111111111010","000000000000001110","111111111111111101","000000000000011010","000000000000010101","111111111111111010","000000000000001001","111111111111111011","000000000000101100","111111111111101101","000000000000001000","111111111111110011","111111111111110110","000000000000000101","000000000000000011","111111111111111101","111111111111101110","000000000000010100","000000000000000010","111111111111100100","111111111111101001","111111111111100101","111111111111100111","000000000000100000","000000000000001110","111111111111110110","000000000000100000","111111111111111001","000000000000100010","111111111111100011","111111111111111011","111111111111111010","000000000000011100","111111111111110100","000000000000000000","000000000000100001","111111111111100011","000000000000000001","111111111111101010","111111111111101111","000000000000001101","111111111111111100","111111111111111101","111111111111100001","000000000000000011","000000000000000111","000000000000000000","111111111111110000","000000000000000010","000000000000011010","111111111111110101","000000000000000101","000000000000101111","000000000001000101","111111111111001110","111111111111110010","111111111111011000","111111111111110001","111111111111101111","000000000000100011","000000000000010110","111111111111110001","111111111111001001","111111111111111000","000000000000010110","111111111111100101","000000000000110000","000000000000010001","000000000000000001","000000000000000010","000000000000000001","111111111111111011","111111111111001110","000000000000000011","000000000001000111","111111111111101101","111111111111101100","000000000000001000","111111111111010100","000000000000010001","000000000000001101","111111111111110101","000000000000001111","111111111111111100","000000000000011110","111111111111110101","111111111111000111","111111111111110100","111111111111011000","111111111111011110","111111111111110011","111111111111100000","111111111111101100","111111111111100011","111111111111110101","000000000000101000","111111111111110000","000000000000011101","000000000000011000","111111111111110111","111111111111010100","111111111111101111","000000000000001100","000000000000010110","111111111111111110","111111111111011100","111111111111110001","111111111111110000","111111111111111001","000000000000010100","111111111111011011","111111111111100101","000000000000011101","000000000000001101","111111111111111110","111111111111111110","111111111111111000","111111111111100111","000000000000001011","000000000000001001","000000000000101001","000000000000001001","000000000000010000","111111111111001110","000000000000001000","111111111111111001"),
("000000000000001101","111111111111101001","111111111111110111","000000000000000011","000000000000000000","000000000000100001","000000000000000000","111111111111101011","000000000000100110","111111111111101111","000000000000001001","111111111111110100","000000000000000101","111111111111101001","111111111111111101","000000000000011000","111111111111111000","111111111111111101","000000000000011100","000000000000001111","000000000000100010","111111111111101111","111111111111111001","111111111111111011","111111111111100001","000000000000101011","000000000000000011","000000000000000111","000000000000000011","111111111111100111","000000000000101011","111111111111110011","111111111111110110","111111111111111100","000000000000100111","111111111111101101","111111111111110111","000000000000101011","111111111111110101","111111111111011000","000000000000000110","111111111111111111","000000000000011110","000000000000011100","000000000000001001","111111111111100110","111111111111111011","000000000000100110","111111111111101000","111111111111111100","000000000000011011","000000000000000110","000000000000000000","000000000000001100","000000000000000101","000000000000010101","111111111111110110","000000000000000001","111111111111101011","000000000000000000","111111111111011111","000000000000000100","000000000000001010","000000000000000111","111111111111110000","000000000000000000","111111111111111011","111111111111101111","000000000000000000","111111111111111100","000000000000100110","111111111111111000","111111111111011001","000000000000001011","111111111111101110","000000000000000101","000000000000001010","000000000000000101","111111111111101011","000000000000011010","111111111111100100","000000000000001110","000000000000010110","111111111111011101","111111111111110000","111111111111110101","111111111111111011","000000000000100000","111111111111100001","111111111111101001","111111111111100011","111111111111111000","111111111111110000","000000000000011010","111111111111101001","111111111111111111","000000000000000110","000000000000011010","111111111111111101","111111111111111010","000000000000011110","111111111111101100","000000000000001001","000000000000010111","000000000000000000","000000000000011101","000000000000000111","000000000000000000","000000000000000010","111111111111110101","000000000000001001","000000000000010100","000000000000001011","000000000000000000","000000000000001110","000000000000100110","000000000000011101","000000000000010000","111111111111110100","111111111111111010","111111111111110111","000000000000101010","000000000000010001","111111111111101111","000000000000001111","000000000000000001","000000000000001011","000000000000001001"),
("111111111111110010","000000000000001000","111111111111111000","111111111111110001","111111111111101111","111111111111101110","000000000000001111","000000000000000010","111111111111111011","000000000000001110","111111111111111011","000000000000001110","111111111111110011","000000000000000101","111111111111110110","111111111111111001","111111111111111110","000000000000011000","111111111111111011","000000000000011001","000000000000001101","000000000000010001","111111111111101110","111111111111110111","111111111111110001","000000000000000000","111111111111111110","000000000000000100","000000000000000110","111111111111110111","000000000000010010","111111111111100110","111111111111110010","000000000000000110","111111111111111000","111111111111111111","000000000000000010","000000000000000001","000000000000000011","111111111111111101","111111111111111010","000000000000000111","111111111111100111","111111111111111111","111111111111111010","000000000000000110","111111111111110011","000000000000001001","000000000000010000","000000000000001110","111111111111111011","000000000000010010","000000000000010100","111111111111101110","111111111111111011","111111111111101110","000000000000010011","000000000000001011","111111111111110110","000000000000001101","111111111111110011","000000000000000011","000000000000000000","000000000000001001","000000000000000101","000000000000001100","111111111111110010","000000000000001010","000000000000001111","111111111111111110","111111111111101011","000000000000010101","111111111111111011","000000000000001000","111111111111111101","111111111111101011","000000000000000101","111111111111110100","000000000000000101","111111111111111001","111111111111110010","000000000000000001","000000000000000111","111111111111110110","000000000000001110","000000000000001101","000000000000000010","111111111111110011","000000000000001000","000000000000000110","000000000000001101","000000000000001110","000000000000001100","000000000000001111","000000000000000000","111111111111101011","111111111111110101","111111111111110001","000000000000011110","111111111111100101","111111111111111110","000000000000010001","111111111111110100","000000000000000000","000000000000010101","111111111111110011","000000000000000000","111111111111111000","111111111111110111","000000000000001110","111111111111111001","111111111111111111","000000000000001111","000000000000001010","000000000000000011","000000000000000111","111111111111111010","000000000000010100","111111111111111101","000000000000010111","000000000000001000","000000000000010111","000000000000000010","000000000000000010","000000000000000111","000000000000000111","000000000000001101","111111111111100101"),
("111111111111110100","111111111111111011","000000000000000110","111111111111111101","111111111111110111","111111111111101011","000000000000000110","111111111111111111","111111111111111011","000000000000000000","111111111111111010","000000000000011000","111111111111111101","000000000000001111","000000000000000000","000000000000000000","000000000000010011","111111111111100101","000000000000000111","000000000000001000","000000000000001001","000000000000001110","111111111111111011","111111111111101110","000000000000010001","111111111111101001","000000000000001001","111111111111100010","000000000000001010","111111111111111111","111111111111111101","111111111111111010","111111111111111101","111111111111110101","000000000000000100","000000000000010100","000000000000010001","000000000000001110","000000000000000000","000000000000011111","000000000000010111","111111111111110100","000000000000010110","000000000000001111","000000000000001100","000000000000001000","000000000000001101","111111111111111010","000000000000001100","000000000000011001","111111111111111101","111111111111111101","000000000000011011","000000000000010000","000000000000000011","111111111111110010","000000000000000110","000000000000001111","000000000000010100","111111111111111111","000000000000011101","111111111111011110","000000000000000101","000000000000000010","111111111111111010","111111111111111011","000000000000001010","000000000000011100","000000000000010110","000000000000000100","000000000000000000","000000000000010010","000000000000011100","000000000000010101","000000000000011011","111111111111110011","111111111111110000","111111111111111010","111111111111111010","000000000000010000","111111111111101011","111111111111111011","111111111111110110","000000000000000001","111111111111110100","000000000000000100","000000000000000010","111111111111110111","000000000000001011","000000000000000101","111111111111110101","000000000000001110","000000000000001100","000000000000000010","111111111111101101","000000000000010110","111111111111111100","000000000000000111","000000000000011101","000000000000011101","111111111111111100","111111111111101010","111111111111111010","111111111111101100","000000000000000100","111111111111101011","000000000000010000","000000000000000111","000000000000010100","111111111111100101","000000000000010000","111111111111101000","000000000000000000","000000000000010110","000000000000010100","111111111111011011","111111111111110100","000000000000011101","000000000000010110","111111111111111111","111111111111111000","111111111111110101","000000000000000000","000000000000010110","000000000000010000","111111111111101001","111111111111100101","000000000000010000"),
("111111111111111110","111111111111010111","111111111111110011","111111111111111010","111111111111110011","111111111111100010","111111111111100100","111111111111001010","000000000000011000","000000000000010111","000000000000010111","111111111111110101","000000000000011100","000000000000100101","000000000000010101","000000000000001011","111111111111100100","000000000000011010","000000000000010100","000000000000011101","000000000000011101","000000000000111110","111111111111111110","000000000000000100","000000000000100011","111111111111110110","111111111111110101","111111111111011111","000000000000000001","111111111111110110","111111111111101111","000000000000110110","111111111111100010","000000000000001010","000000000000010001","111111111111110011","000000000000000011","111111111111111010","111111111111110101","000000000000100011","000000000000100101","000000000000100011","000000000000100100","000000000000010011","111111111111101001","000000000000010001","111111111111111101","000000000000001100","000000000000001101","000000000000100001","000000000000000011","111111111111101010","000000000000101101","000000000000001000","000000000000001000","000000000000000100","111111111111101010","000000000000011111","000000000000001101","111111111111110110","000000000000010111","111111111111110111","111111111111110101","111111111111111001","000000000000011011","000000000000011001","111111111111101011","111111111111011111","111111111111111100","000000000000000110","111111111111010111","000000000000000000","000000000000001010","000000000000001011","111111111111110110","111111111111110000","111111111111101011","111111111111110000","000000000000010011","000000000000001011","000000000000000001","111111111111101001","111111111111100111","000000000000100001","111111111111010000","000000000000001100","000000000000001010","111111111111110111","111111111111100100","000000000000001111","000000000000011100","111111111111110000","000000000000010001","000000000000001000","111111111111110001","111111111111111011","111111111111100110","111111111111100111","000000000000001001","000000000000111001","111111111111111011","111111111111101101","111111111111110101","111111111111001111","000000000000001001","111111111111101111","111111111111101111","000000000000010100","111111111111111000","000000000000010101","111111111111110100","111111111111011010","111111111111100001","000000000000010101","111111111111111111","111111111111011111","111111111111011001","000000000000000010","000000000000000000","000000000000100001","000000000000010001","111111111111110010","111111111111111110","000000000000111011","000000000000011111","111111111111101101","000000000000001000","111111111111110101"),
("111111111111110011","111111111111100011","000000000000000100","000000000000001110","000000000000000000","000000000000010100","000000000000000101","000000000000000111","111111111111100110","000000000000100001","111111111111100000","111111111111101101","000000000000000101","000000000000100010","000000000000001101","111111111111111001","000000000000001001","000000000000001000","111111111111111000","000000000000001011","000000000000010001","000000000000000110","111111111111100101","111111111111100110","000000000000001011","000000000000001110","000000000000010111","000000000000000110","000000000000001001","000000000000010010","000000000000011101","000000000000100011","111111111111110011","111111111111100001","000000000000000111","111111111111100111","000000000000000101","111111111111101101","111111111111011100","111111111111111101","111111111111110011","111111111111111101","000000000000010001","111111111111111101","111111111111111100","000000000000010110","111111111111100010","000000000000000111","111111111111111010","000000000000001001","111111111111101011","111111111111101010","111111111111110010","000000000000001001","000000000000100001","000000000000001010","111111111111100110","000000000000001001","111111111111101111","000000000000000000","000000000000000101","000000000000001011","000000000000000110","000000000000000110","111111111111110110","111111111111110001","000000000000001010","111111111111100001","111111111110111100","000000000000001010","000000000000010011","111111111111101111","000000000000011101","000000000000100001","111111111111111001","111111111111100111","000000000000001001","111111111111101101","111111111111101011","111111111111100101","111111111111101110","111111111111110001","000000000000011001","000000000000011100","111111111111111111","000000000000001111","000000000000011011","000000000000010001","111111111111110000","000000000000100001","000000000000000000","111111111111101110","111111111111111011","111111111111100101","000000000000010110","111111111111100001","000000000000001110","111111111111111001","000000000000010011","000000000000000110","111111111111111010","111111111111011001","111111111111011110","111111111111111001","111111111111111011","111111111111101000","000000000000001100","111111111111100101","111111111111100110","111111111111100011","000000000000010101","000000000000011010","111111111111101110","111111111111111111","000000000000001100","111111111111110111","111111111111110010","000000000000010001","111111111111110110","111111111111111101","111111111111110100","111111111111111010","000000000000001110","000000000000001111","000000000000100101","111111111111101110","111111111111111100","000000000000000101"),
("000000000000000111","000000000000100000","000000000000001100","111111111111111011","000000000000101001","000000000000000100","111111111111111100","000000000000011110","111111111111100101","000000000000000001","111111111111110010","111111111111110010","111111111110110101","000000000000000011","000000000000010101","111111111111110101","111111111111111011","111111111111101111","000000000000000000","111111111111101010","111111111111101010","000000000000000100","000000000000010010","111111111111011111","111111111111111100","111111111111101101","000000000000010111","111111111111101110","000000000000000000","000000000000011010","111111111111111110","111111111111101110","111111111111110011","000000000000000100","111111111111010101","111111111111100001","111111111111111100","111111111111110100","000000000000000010","000000000000000000","000000000000010010","000000000000011001","000000000000001000","111111111111010011","111111111111111010","000000000000001101","111111111111101001","111111111111101110","000000000000001011","000000000000000000","111111111111000110","000000000000001111","111111111111111110","000000000000000000","000000000000000110","000000000000011001","111111111111101101","111111111111100011","000000000000010000","111111111111110000","111111111111110111","000000000000001000","000000000000001100","111111111111111111","111111111111111000","000000000000100010","111111111111101110","111111111111001001","111111111110110111","000000000000000001","111111111111011110","111111111111101110","000000000000000000","000000000000010001","111111111111100010","111111111111011010","111111111111110111","111111111111110101","111111111111111001","111111111111101110","111111111111111100","000000000000010010","111111111111111100","000000000000011100","111111111111111010","111111111111101111","000000000000010010","000000000000001010","111111111111001110","111111111111111011","111111111111111110","000000000000000110","000000000000000001","000000000000001011","000000000000010110","000000000000000010","111111111111101111","111111111111110010","111111111111111101","000000000000001110","000000000000010101","111111111111100110","111111111111111111","111111111111101101","111111111111010101","111111111111101010","000000000000000000","111111111111111011","000000000000000110","111111111111110001","000000000000011010","000000000000101110","111111111111111010","000000000000001010","111111111111100111","000000000000001110","111111111111101011","111111111111111000","111111111111100010","111111111111101111","111111111111100111","000000000000000110","000000000000001111","111111111111110011","111111111111101011","000000000000000000","111111111111110010","000000000000000000"),
("000000000000000110","000000000000010101","000000000000010011","111111111111110000","000000000000010100","000000000000000100","111111111111111010","000000000000000100","111111111111000100","000000000000100000","111111111110111011","000000000000000110","111111111111000101","111111111111100011","000000000000001001","111111111111011010","000000000000001100","111111111111101001","111111111111110011","000000000000000101","000000000000000100","000000000000001000","000000000000011110","111111111111111001","000000000000011010","111111111111100000","000000000000001101","111111111111101010","000000000000000000","111111111111101110","111111111111011101","111111111111110010","111111111111101101","111111111111010001","111111111111100110","111111111111111001","000000000000000110","111111111111010001","111111111111110001","000000000000000010","111111111111110010","111111111111110011","111111111111110110","111111111111000111","000000000000010101","111111111111111010","000000000000000100","000000000000011011","000000000000010001","000000000000000101","000000000000001101","000000000000010111","111111111111111010","111111111111101110","111111111111010001","000000000000000111","111111111111011011","000000000000001100","000000000000100100","000000000000001100","000000000000000011","000000000000101011","111111111111101110","111111111111110111","111111111111001111","000000000000011001","111111111111111010","111111111111110100","111111111110010001","000000000000000011","111111111111101101","111111111111010000","000000000000110010","111111111111101101","111111111111110010","111111111111110011","000000000000000000","111111111111111111","000000000000010000","000000000000011100","111111111111111010","000000000000000101","111111111111111011","111111111111011001","111111111111111000","111111111111111000","000000000000011000","111111111111110101","111111111111001110","000000000000001110","000000000000010010","111111111111100100","111111111111111110","000000000000100111","111111111111110101","111111111111101111","000000000000000101","111111111111110011","111111111111011001","111111111111111110","000000000000001000","000000000000100011","111111111111111011","111111111111110101","111111111111100110","000000000000001101","000000000000001101","111111111111110010","111111111111111100","111111111111111001","000000000000000110","000000000000000000","000000000000000101","000000000000001010","111111111111101011","000000000000100011","111111111111110011","111111111111101010","111111111111100001","111111111111010110","111111111111011101","111111111111111100","111111111111111111","000000000000010110","111111111111110011","111111111111111000","111111111111010001","111111111111111100"),
("000000000000101100","000000000000110001","000000000000100110","111111111111111111","000000000000001100","000000000000010011","000000000000001010","000000000000011100","111111111111010001","000000000000111100","111111111111001101","000000000000010110","111111111111101110","000000000000010100","000000000000011010","000000000000000000","000000000000001000","000000000000001010","111111111111101010","111111111111100101","000000000000000011","000000000000000101","000000000000000101","111111111111100000","111111111111111101","000000000000001010","000000000000001100","000000000000000001","111111111111100001","111111111111111100","000000000000000111","000000000000000110","111111111111110000","111111111111100000","111111111111111110","111111111111101101","111111111111101011","111111111111111000","111111111111101001","000000000000000000","111111111111110000","000000000000001000","111111111111100010","111111111111000110","000000000000000101","000000000000010000","111111111111100111","000000000000101000","111111111111101101","111111111111101011","000000000000011001","000000000000011101","000000000000001011","111111111111011011","111111111111000011","111111111111101100","111111111111100001","111111111111101011","000000000000001010","111111111111111101","111111111111101110","000000000001001000","111111111111101001","000000000000010100","111111111110111101","111111111111111100","000000000000011111","000000000000010000","111111111110100111","000000000000011111","000000000000010111","111111111111011111","000000000000011100","000000000000000001","111111111111111010","000000000000001001","111111111111111001","000000000000001000","111111111111110000","000000000000001100","000000000000000011","000000000000000011","000000000000011001","111111111111001000","000000000000000011","111111111111111110","000000000000101100","111111111111111011","111111111111111000","111111111111110011","111111111111110011","111111111111101001","000000000000000000","111111111111111111","000000000000010010","111111111111011110","000000000000010010","000000000000000110","111111111111101000","111111111111110000","000000000000101001","000000000000001100","111111111111100111","000000000000001010","111111111111010110","000000000000010100","000000000000010111","000000000000000101","000000000000000000","000000000000000111","000000000000001111","111111111111110110","111111111111111111","111111111111110111","111111111111110101","111111111111111110","111111111111111001","111111111111101001","111111111111100111","111111111111101001","111111111111001110","111111111111111001","111111111111100110","000000000000001111","000000000000000100","111111111111111000","111111111111100111","000000000000000111"),
("000000000000000111","000000000000110000","000000000000110110","111111111111110010","000000000000000110","000000000000000101","000000000000001100","000000000000001110","111111111111001101","000000000000101011","111111111110110000","000000000000011110","111111111111110110","000000000000001100","000000000000000001","000000000000000100","111111111111111000","000000000000001000","111111111111101010","111111111111110100","111111111111110011","000000000000010011","000000000000001001","111111111111101010","000000000000011010","111111111111110101","000000000000010100","111111111111111110","111111111111110110","000000000000000000","111111111111110111","111111111111101010","111111111111110011","111111111111110000","111111111111101110","111111111111111111","111111111111111101","111111111111111011","111111111111100101","000000000000000010","111111111111111011","111111111111111110","111111111111001110","111111111111010101","000000000000001101","111111111111111000","111111111111011011","000000000000010011","111111111111110110","111111111111101000","111111111111111111","000000000000011010","000000000000010011","111111111111011011","111111111111110011","111111111111111111","111111111111101111","000000000000000111","000000000000011010","000000000000000000","000000000000000000","000000000000101001","000000000000001011","000000000000010101","111111111111101100","000000000000011110","000000000000010011","000000000000010100","111111111110111100","000000000000000111","000000000000001010","111111111111101011","000000000000000110","111111111111110110","111111111111100111","000000000000100011","000000000000000100","111111111111110101","000000000000001100","111111111111111110","000000000000011001","111111111111111101","000000000000110001","111111111111011101","000000000000000100","000000000000011000","000000000000011110","000000000000001101","111111111111110111","111111111111101001","111111111111110101","000000000000001100","000000000000000101","000000000000011110","000000000000000110","111111111111100110","111111111111111011","111111111111111010","111111111111000011","000000000000001000","000000000000101000","000000000000010101","111111111111110001","000000000000010000","111111111111010010","000000000000000001","000000000000010000","000000000000001011","000000000000011001","000000000000010110","000000000000000101","000000000000001001","111111111111110110","111111111111100001","111111111111101111","111111111111111001","111111111111101111","111111111111110011","111111111111101110","111111111111100100","111111111111110111","111111111111111101","111111111111101101","111111111111111011","000000000000001110","000000000000010000","111111111111100111","111111111111111101"),
("000000000000001111","000000000000100000","000000000000101111","000000000000000011","000000000000011011","000000000000001100","000000000000011011","000000000000001001","111111111111011101","000000000000111101","111111111110011111","000000000000011100","111111111111101111","000000000000010101","000000000000001110","111111111111111011","000000000000000101","111111111111110111","111111111111100110","111111111111111000","111111111111110100","000000000000111001","000000000000001011","111111111111101111","111111111111111110","000000000000000010","000000000000010000","111111111111110000","000000000000000010","000000000000011011","111111111111111110","111111111111100011","111111111111101010","000000000000000000","111111111111111011","111111111111110101","111111111111110001","000000000000000000","000000000000010111","000000000000001001","111111111111100001","111111111111111110","111111111111010100","111111111111101111","111111111111111110","000000000000000100","111111111111010011","000000000000001011","111111111111111110","111111111111111101","000000000000011000","000000000000010001","000000000000010110","111111111111100111","111111111111110011","000000000000000000","111111111111110010","000000000000000110","000000000000010111","000000000000010001","000000000000000010","000000000000001110","000000000000010111","000000000000010110","111111111111110001","000000000000011010","000000000000010000","000000000000000101","111111111111011000","111111111111111111","000000000000000101","111111111111110000","111111111111111011","111111111111111101","000000000000001011","000000000000010101","000000000000000000","111111111111110100","000000000000010111","000000000000010101","000000000000011010","111111111111111010","000000000000100100","111111111111101001","000000000000001011","000000000000010101","000000000000010110","000000000000000011","000000000000001100","000000000000100001","000000000000011011","000000000000000000","000000000000010010","000000000000001001","000000000000000000","000000000000001001","111111111111101101","111111111111111001","111111111111011001","000000000000000000","000000000000010010","000000000000101100","000000000000001001","000000000000000000","111111111111101111","000000000000001001","000000000000010111","111111111111100101","000000000000011100","000000000000010001","111111111111110111","111111111111101001","000000000000001110","111111111111101111","000000000000000101","000000000000000000","111111111111101001","111111111111010111","000000000000000111","000000000000000000","111111111111110000","111111111111100110","111111111111110001","000000000000011010","000000000000001110","111111111111111010","111111111111110000","000000000000001101"),
("000000000000010011","111111111111110001","000000000000100101","111111111111101011","000000000000000010","111111111111111010","000000000000010101","111111111111101011","111111111111100111","000000000000001110","111111111110000110","000000000000010100","111111111111010011","000000000000011010","000000000000001101","111111111111110010","000000000000101100","111111111111100101","111111111111011011","000000000000001111","111111111111110001","000000000000101001","000000000000001010","111111111111111010","000000000000001100","000000000000000010","000000000000010101","111111111111111010","111111111111111101","000000000000100110","111111111111111100","000000000000000010","111111111111011100","000000000000001011","111111111111110001","000000000000000010","111111111111110101","111111111111011011","000000000000100111","111111111111101100","000000000000000101","111111111111101000","111111111111011000","111111111111101100","111111111111110101","000000000000010000","111111111111011011","000000000000001111","000000000000011010","000000000000001010","000000000000010010","000000000000001000","000000000000010001","111111111111100011","111111111111110010","111111111111110100","000000000000100010","000000000000000100","000000000000001101","000000000000010001","111111111111101010","000000000000100111","000000000000100101","000000000000001011","000000000000001100","000000000000010010","000000000000000001","000000000000011110","000000000000001011","000000000000010000","111111111111110001","111111111111100111","000000000000010001","111111111111110010","111111111111110001","111111111111111111","000000000000000011","000000000000000000","000000000000000101","000000000000001001","000000000000101000","111111111111101110","000000000000011001","111111111111011111","000000000000000100","000000000000011000","000000000000100101","000000000000011110","000000000000010110","000000000000011001","000000000000101100","111111111111101101","000000000000100011","000000000000011001","000000000000001010","111111111111101111","111111111111100100","111111111111111110","000000000000011011","000000000000001001","000000000000101101","000000000000010101","000000000000001010","111111111111101101","111111111111110111","111111111111111001","111111111111111100","111111111111111101","000000000000011000","000000000000001110","111111111111111000","111111111111101100","111111111111111110","111111111111100000","000000000000010011","000000000000011111","111111111111110010","111111111111100101","000000000000010010","000000000000001101","111111111111001110","111111111111101110","000000000000000100","000000000000001010","000000000000010000","000000000000000110","111111111111011111","000000000000000001"),
("111111111111110111","111111111111010010","000000000000011111","000000000000000000","000000000000001111","111111111111110100","000000000000010111","111111111111010111","111111111111100001","000000000000010111","111111111110101000","000000000000011000","111111111111001111","111111111111110011","000000000000001101","000000000000011000","000000000000101000","111111111111111001","111111111111010011","000000000000001000","111111111111111010","111111111111111100","111111111111100110","111111111111100011","000000000000010011","111111111111101100","000000000000001011","111111111111011110","000000000000001110","000000000000000111","000000000000000110","111111111111101011","000000000000000011","000000000000100010","111111111111111011","111111111111101110","000000000000001010","111111111111101111","000000000000011101","111111111111111110","000000000000001011","111111111111101010","000000000000000111","000000000000001010","000000000000000101","000000000000100010","111111111111011100","000000000000010101","000000000000011001","000000000000000101","000000000000111000","000000000000000101","000000000000100010","111111111111101001","111111111111111010","111111111111101111","000000000000010010","000000000000000111","111111111111111111","000000000000000101","111111111111111000","000000000000011101","000000000000010110","000000000000000101","000000000000000101","000000000000010010","000000000000000100","000000000000011110","000000000000010100","000000000000010010","111111111111101001","111111111111010101","111111111111101110","111111111111110100","000000000000000000","000000000000010001","000000000000010001","111111111111101110","000000000000000010","111111111111110010","111111111111111101","111111111111110001","000000000000001001","111111111111001111","111111111111011110","000000000000011001","000000000000000100","000000000000010001","000000000000100100","000000000000001111","000000000000010001","111111111111110101","000000000000011001","000000000000001011","000000000000000011","111111111111100111","111111111111010101","111111111111111100","000000000000010000","111111111111110110","000000000000111000","000000000000001001","111111111111110101","000000000000000000","000000000000000100","000000000000011001","000000000000000010","111111111111110110","000000000000011011","000000000000010110","111111111111110010","111111111111000101","000000000000001010","000000000000000110","111111111111110111","000000000000000011","111111111111111110","111111111111111011","000000000000011101","000000000000000110","111111111111100001","000000000000000101","000000000000010101","000000000000000011","000000000000110001","000000000000010001","111111111111111001","000000000000000000"),
("111111111111101111","111111111110111110","000000000000000110","000000000000001000","111111111111111111","000000000000011001","000000000000001010","111111111111100001","111111111111101011","111111111111100111","111111111110100011","000000000000001000","111111111111001100","111111111111110011","000000000000000110","000000000000001101","000000000000110001","111111111111111111","111111111111001101","000000000000000011","000000000000000010","111111111111100000","111111111111101011","000000000000001100","000000000000001100","111111111111110010","000000000000000000","111111111111110011","111111111111110010","000000000000100010","000000000000000011","111111111111101101","111111111111111111","000000000000011100","000000000000000101","000000000000000011","000000000000000010","111111111111111010","000000000000010110","111111111111110000","111111111111011100","111111111111110111","111111111111111001","111111111111111100","000000000000010101","111111111111111100","000000000000000001","000000000000100011","000000000000010000","000000000000011011","000000000000011101","000000000000010001","000000000000000111","111111111111111010","111111111111111001","000000000000000001","000000000000000111","111111111111100100","000000000000011100","111111111111111111","111111111111111100","000000000000001111","000000000000110011","000000000000011101","000000000000010111","000000000000001011","111111111111110000","000000000000011110","000000000000011000","000000000000010011","111111111111111001","111111111111100110","111111111111111010","111111111111110100","111111111111100100","000000000000100011","000000000000011000","111111111111110100","000000000000000100","000000000000000010","111111111111111011","000000000000011011","111111111111111001","000000000000001110","000000000000000101","111111111111110010","000000000000011100","111111111111101000","000000000000001111","000000000000010011","000000000000000100","111111111111110110","000000000000001011","111111111111111101","111111111111111110","111111111111101000","111111111111101010","000000000000011111","000000000000100111","111111111111111111","000000000000010011","000000000000011011","111111111111111010","000000000000000111","000000000000000011","000000000000000101","000000000000010110","111111111111111110","000000000000001000","000000000000011000","000000000000010001","111111111111100101","000000000000000110","000000000000000110","000000000000010010","000000000000101010","000000000000001110","111111111111011100","000000000000011011","111111111111110001","111111111111101001","000000000000000110","111111111111100110","111111111111000110","000000000000110000","000000000000100011","000000000000010111","111111111111101111"),
("000000000000010001","111111111111000011","111111111111110011","111111111111111101","111111111111111101","000000000000000010","000000000000010011","111111111111111101","000000000000000110","111111111111100101","111111111111011000","000000000000001100","111111111111000111","111111111111101110","111111111111010110","000000000000101010","000000000000111011","111111111111111101","111111111111100110","111111111111110001","111111111111111010","111111111111100101","111111111111001011","000000000000000111","111111111111111000","000000000000000101","000000000000010110","111111111111100011","111111111111111000","000000000000001111","000000000000000101","111111111111111011","000000000000100001","111111111111110000","111111111111111101","000000000000100111","000000000000001001","000000000000001011","000000000000000111","000000000000001011","111111111111110010","111111111111101000","000000000000010100","000000000000000000","000000000000100000","111111111111110001","000000000000110010","000000000000011100","111111111111111101","000000000000101010","000000000000001100","000000000000010100","000000000000000100","111111111111110101","111111111111101111","111111111111101110","000000000000010000","111111111111110001","000000000000010011","000000000000001110","111111111111111111","000000000000001000","000000000000100000","000000000000011100","000000000000011011","000000000000000010","000000000000000001","000000000000001111","000000000000110101","111111111111100010","000000000000010100","111111111111011001","000000000000010100","111111111111111111","000000000000000000","000000000000011111","000000000000010000","000000000000000001","000000000000000000","000000000000000011","111111111111111011","000000000000010100","000000000000000010","000000000000011010","111111111111111011","000000000000001101","000000000000011111","000000000000001111","111111111111110000","000000000000011001","111111111111101101","000000000000001111","000000000000000000","000000000000001011","111111111111101100","111111111111111101","111111111111110011","111111111111111010","000000000000101101","111111111111111111","000000000000010010","000000000000010101","000000000000001000","000000000000000001","111111111111111101","000000000000100110","000000000000001011","111111111111101101","000000000000011001","000000000000000110","111111111111111111","111111111111001101","000000000000010100","000000000000001000","000000000000010100","000000000000000100","111111111111111100","111111111111011101","000000000000101001","000000000000000010","111111111111101011","000000000000011011","111111111111101100","111111111110011001","000000000000101000","111111111111111011","000000000000001110","000000000000001110"),
("000000000000011001","111111111111101001","111111111111100010","000000000000010100","111111111111101101","000000000000011011","000000000000000011","111111111111101011","000000000000010000","111111111111011110","000000000000001100","111111111111110001","111111111111101100","000000000000010011","111111111111100100","000000000000001101","111111111111111010","000000000000011000","111111111111101010","000000000000000111","111111111111110110","111111111111100100","111111111110111101","000000000000001011","000000000000001010","000000000000011110","000000000000000111","000000000000000111","000000000000010110","111111111111111000","000000000000001111","000000000000000000","000000000000000011","111111111111100110","111111111111101011","000000000000110100","111111111111101111","000000000000011000","000000000000010110","111111111111110100","111111111111011010","000000000000000010","000000000000010010","000000000000000011","000000000000001110","111111111111100001","000000000000111011","000000000000101101","111111111111110000","000000000000100111","111111111111011010","000000000000001110","111111111111100011","000000000000000000","000000000000001011","000000000000010000","000000000000011111","000000000000010000","111111111111111001","111111111111101010","111111111111111001","000000000000010011","111111111111110110","000000000000010110","000000000000100101","000000000000000010","000000000000000000","000000000000010111","000000000000100010","111111111111010010","000000000000010000","111111111111111101","000000000000000000","000000000000000101","000000000000000011","000000000000001100","000000000000001100","000000000000001011","111111111111111010","111111111111110101","000000000000001101","111111111111111001","000000000000000111","000000000000110110","000000000000100001","111111111111111000","000000000000010010","111111111111110001","111111111111110101","000000000000001101","111111111111110000","000000000000100101","111111111111110101","000000000000000000","000000000000001000","000000000000100111","111111111111101100","000000000000001101","000000000000000110","000000000000001000","000000000000001000","000000000000000100","000000000000011010","000000000000010010","000000000000011011","000000000000000011","000000000000010111","111111111111101110","000000000000001010","000000000000000100","000000000000001110","111111111111110001","000000000000000111","000000000000001101","000000000000001001","000000000000001100","000000000000011101","111111111111101111","000000000000101111","111111111111110110","111111111111100011","000000000000001010","000000000000000001","111111111110010011","000000000000011001","111111111111100100","000000000000010000","111111111111110111"),
("000000000000011110","111111111111111100","111111111111101000","000000000000000011","111111111111101000","000000000000000110","111111111111110101","000000000000010100","000000000000100100","111111111111110010","111111111111110100","111111111111111110","111111111111111111","000000000000010101","111111111111101011","000000000000000100","111111111111111111","000000000000001111","111111111111111111","111111111111101001","111111111111101111","111111111111110101","111111111110111111","000000000000011111","111111111111111011","000000000000011010","000000000000011001","000000000000010000","000000000000011101","111111111111111101","000000000000000001","000000000000001000","000000000000001001","111111111111110011","000000000000100100","000000000000101111","111111111111111110","000000000000101011","000000000000010001","000000000000001000","111111111111110110","000000000000110001","000000000000010011","000000000000000111","000000000000010100","000000000000000010","000000000000110011","000000000000010000","000000000000000000","111111111111111100","111111111111101101","000000000000010101","111111111111011001","000000000000000001","000000000000011100","000000000000011100","000000000000010110","111111111111111010","111111111111100010","111111111111101010","111111111111111101","000000000000011110","111111111111101011","000000000000010000","000000000000110000","111111111111111011","000000000000010000","000000000000011101","000000000000011100","111111111111010010","000000000000011110","000000000000011110","111111111111111011","000000000000010001","000000000000010001","000000000000010001","000000000000010100","111111111111111111","000000000000001001","000000000000001001","111111111111111011","000000000000010010","111111111111110100","000000000000100101","000000000000010101","111111111111111010","000000000000010011","000000000000001010","000000000000000101","000000000000001001","111111111111101110","000000000000000000","111111111111100000","111111111111101000","000000000000000000","000000000000000111","000000000000000100","000000000000010110","111111111111110000","000000000000101110","000000000000000100","000000000000000010","111111111111111101","000000000000101000","000000000000011110","111111111111111101","000000000000010010","000000000000011101","000000000000110001","111111111111100001","111111111111111011","111111111111100111","000000000000011001","000000000000010111","000000000000001000","000000000000100010","000000000000001001","000000000000000111","000000000000011001","000000000000010111","000000000000000010","111111111111111010","000000000000100010","111111111111010001","000000000000001100","111111111111101110","000000000000010001","111111111111111100"),
("000000000000011011","111111111111110000","000000000000000000","000000000000000111","000000000000001010","000000000000011010","000000000000011000","000000000000010001","000000000000001101","111111111111110101","111111111111111000","111111111111111110","000000000000000110","000000000000001001","000000000000010100","111111111111100000","111111111111100001","000000000000001111","000000000000010000","111111111111100100","000000000000000011","000000000000000000","111111111111100101","000000000000100011","111111111111110101","000000000000101001","000000000000001101","000000000000011101","000000000000001000","111111111111111111","000000000000000110","000000000000010110","111111111111111000","000000000000001111","000000000000000001","000000000000100100","111111111111110000","000000000000001110","000000000000010001","000000000000011010","111111111111111001","000000000000001000","000000000000000010","000000000000000111","000000000000001100","000000000000011000","000000000000001111","000000000000010001","111111111111110111","000000000000011000","000000000000001000","000000000000000001","111111111111110010","000000000000001100","000000000000010000","000000000000010010","000000000000011001","111111111111111000","111111111111100000","111111111111101010","000000000000001100","000000000000000111","111111111111100010","111111111111111001","000000000000100010","111111111111111101","000000000000000100","111111111111110111","000000000000011000","111111111111110011","000000000000000100","000000000000000100","111111111111110111","000000000000010000","000000000000010101","111111111111110001","000000000000010000","000000000000001011","000000000000010001","000000000000010010","000000000000000001","000000000000000111","000000000000000000","000000000000101100","111111111111111110","000000000000010011","111111111111110110","000000000000010100","000000000000010101","111111111111110111","000000000000011011","000000000000010110","111111111111111000","111111111111011010","111111111111110100","000000000000011010","111111111111100110","000000000000101110","111111111111111110","000000000000001111","000000000000001110","111111111111110001","111111111111110001","000000000000011001","000000000000000000","111111111111110001","000000000000010010","000000000000010001","000000000000010011","111111111111111010","000000000000001011","111111111111011011","000000000000100000","000000000000010000","111111111111111110","111111111111111000","000000000000010010","111111111111101000","000000000000100000","111111111111110111","000000000000000000","000000000000001001","000000000000101001","000000000000000110","000000000000010110","000000000000000000","111111111111110101","000000000000000100"),
("000000000000011111","111111111111110111","000000000000001101","111111111111111010","000000000000010010","000000000000001001","111111111111111000","000000000000010101","000000000000011010","111111111111110001","111111111111100000","111111111111100110","000000000000000111","000000000000011011","000000000000011011","111111111111101001","111111111111111000","111111111111111011","111111111111111110","111111111111101001","111111111111110110","111111111111010101","111111111111101001","000000000000010101","111111111111101000","000000000000010010","000000000000001011","000000000000011000","000000000000010101","111111111111011001","111111111111111110","000000000000001100","111111111111111110","000000000000001100","000000000000010110","000000000000010011","000000000000001011","111111111111111001","000000000000011110","000000000000001111","111111111111101000","111111111111101111","000000000000001110","000000000000010100","000000000000000111","000000000000011111","111111111111101011","000000000000100111","000000000000000110","000000000000000101","111111111111111001","111111111111110101","111111111111101101","111111111111110101","000000000000010100","000000000000001110","111111111111111111","111111111111100010","111111111111011011","000000000000001111","000000000000000000","000000000000000101","111111111111111101","111111111111111000","000000000000101110","111111111111110010","111111111111111000","111111111111111111","000000000000011110","111111111111110010","000000000000011001","111111111111110010","111111111111101111","000000000000010110","000000000000001000","111111111111110100","000000000000000011","000000000000001010","000000000000100011","000000000000001110","000000000000010001","000000000000000101","000000000000001011","000000000000011000","111111111111101011","000000000000100111","000000000000001011","000000000000010100","000000000000010100","111111111111101011","000000000000011011","111111111111100101","111111111111111000","111111111111010111","000000000000000011","000000000000001000","111111111111111100","000000000000110010","111111111111100000","000000000000001110","000000000000011110","111111111111110001","111111111111101110","111111111111111001","111111111111110000","111111111111111101","000000000000011010","000000000000001001","000000000000010000","111111111111111111","000000000000010001","111111111111100101","000000000000010101","000000000000000000","111111111111111110","000000000000000100","111111111111110000","111111111111101000","000000000000001011","111111111111101110","000000000000000001","000000000000000111","000000000000011000","111111111111111001","000000000000001011","000000000000001110","111111111111111000","000000000000011111"),
("111111111111111110","111111111111111111","000000000000000011","000000000000000100","000000000000000001","000000000000011000","111111111111111111","000000000000001000","000000000000100000","111111111111111000","111111111111011101","111111111111111000","000000000000001100","000000000000000110","000000000000011001","111111111111010001","000000000000010000","111111111111111010","111111111111111011","111111111111110001","111111111111110101","111111111111111010","000000000000000011","111111111111101011","111111111111110100","000000000000000011","000000000000010000","111111111111110010","000000000000000110","111111111111111010","111111111111111110","111111111111110111","000000000000001001","000000000000010010","111111111111110011","111111111111101101","111111111111110110","000000000000000110","000000000000000010","000000000000000000","000000000000000010","111111111111010110","111111111111111101","111111111111110110","000000000000010011","000000000000000100","111111111111110100","000000000000011101","000000000000011100","000000000000000000","111111111111111111","111111111111110001","111111111111110100","111111111111110100","000000000000001011","000000000000110000","111111111111111010","000000000000001010","000000000000001010","111111111111110010","000000000000000000","000000000000010001","111111111111111010","000000000000100010","000000000000010100","000000000000001011","111111111111111011","111111111111101010","000000000000011001","111111111111101101","000000000000001000","000000000000000000","111111111111010111","000000000000011001","000000000000001110","111111111111110110","000000000000010000","000000000000001010","000000000000001100","000000000000001011","000000000000010101","000000000000001111","000000000000001001","000000000000101110","111111111111101001","000000000000110111","000000000000000110","000000000000000111","000000000000000101","111111111111100010","000000000000010101","111111111111111110","111111111111101101","111111111111111110","000000000000001100","000000000000010000","000000000000000000","000000000000011010","111111111111111111","000000000000100000","000000000000001101","000000000000000100","000000000000001000","111111111111101001","111111111111111100","111111111111110011","000000000000101010","000000000000000100","000000000000010110","000000000000011110","000000000000010011","111111111110111101","000000000000010100","000000000000000010","000000000000001111","111111111111111101","111111111111100110","000000000000000000","000000000000001111","000000000000000101","111111111111110001","111111111111110001","000000000000011110","000000000000000110","000000000000011101","111111111111110101","111111111111100111","000000000000010000"),
("000000000000000000","111111111111111111","000000000000001011","000000000000000000","111111111111110010","000000000000001011","000000000000011101","111111111111100111","111111111111101110","111111111111111110","111111111111100011","000000000000000001","000000000000100001","000000000000101011","000000000000100110","111111111111100111","111111111111111011","111111111111110000","111111111111101111","111111111111101100","000000000000000100","111111111111111111","111111111111111010","111111111111110101","111111111111101110","111111111111100101","000000000000000000","000000000000000110","111111111111101110","111111111111101010","111111111111011111","111111111111110001","000000000000100010","000000000000010101","111111111111101110","111111111111010100","111111111111110111","111111111111100000","111111111111111110","000000000000010111","111111111111111000","111111111111110010","000000000000000110","000000000000001111","000000000000011010","111111111111111010","000000000000001111","000000000000001101","000000000000001101","111111111111111111","000000000000010101","111111111111111001","000000000000001011","111111111111111111","111111111111110111","000000000000011111","111111111111110000","000000000000001100","000000000000011101","000000000000000011","111111111111110010","111111111111111010","111111111111111001","000000000000010111","111111111111011101","000000000000011011","111111111111011111","111111111111111000","111111111111110100","111111111111101010","000000000000000000","111111111111101110","111111111111100001","000000000000001111","111111111111111101","111111111111111000","000000000000001001","000000000000001010","000000000000000011","000000000000001110","111111111111101000","000000000000000010","000000000000011110","000000000000011110","000000000000000101","000000000001000010","000000000000001010","000000000000000000","000000000000011100","000000000000001000","111111111111111111","111111111111100110","111111111111100001","000000000000000101","000000000000100101","000000000000001000","111111111111110011","000000000000010001","000000000000011010","111111111111110101","000000000000000101","000000000000010001","111111111111110010","111111111111110000","111111111111101101","000000000000001100","000000000000010100","000000000000010011","000000000000000011","000000000000110000","000000000000011001","111111111111011100","000000000000000110","111111111111110000","111111111111111111","000000000000010001","000000000000010001","000000000000010100","111111111111101010","000000000000001011","111111111111110110","111111111111110001","000000000000000000","111111111111111010","000000000000011010","000000000000011100","111111111111101000","000000000000000111"),
("111111111111100101","000000000000000010","000000000000010000","111111111111101000","000000000000011010","000000000000000111","000000000000001100","111111111111100001","111111111111101001","000000000000001000","111111111111101011","111111111111100111","111111111111110101","000000000000000010","000000000000100000","111111111111101001","000000000000011110","111111111111100010","000000000000000000","111111111111111111","111111111111100111","000000000000000000","111111111111100001","000000000000000101","111111111111111111","111111111111100100","111111111111111011","000000000000001010","111111111111111010","111111111111010111","111111111111101010","000000000000000010","000000000000010110","000000000000010010","111111111111100101","111111111111011000","000000000000001010","111111111111101111","000000000000000001","000000000000000000","111111111111110101","000000000000010000","000000000000010000","111111111111111101","111111111111110111","000000000000000000","000000000000101000","111111111111111010","000000000000100000","000000000000000101","000000000000001101","111111111111110111","000000000000001000","000000000000000000","111111111111101000","000000000000011010","000000000000001000","111111111111111000","000000000000010101","111111111111111010","000000000000010101","111111111111110110","111111111111110100","000000000000000001","111111111110101001","000000000000011001","111111111111100000","111111111111101110","000000000000001010","111111111111100110","000000000000000110","111111111111111010","111111111111101110","111111111111111110","111111111111111101","111111111111111111","111111111111111101","111111111111110010","000000000000001100","111111111111111111","000000000000000000","000000000000001111","000000000000011011","000000000000110110","111111111111101111","000000000000101101","000000000000010101","111111111111111011","000000000000000100","000000000000001100","111111111111100100","111111111111101000","111111111111101100","111111111111111011","000000000000011000","111111111111101101","111111111111110101","000000000000110001","000000000000011001","000000000000010001","111111111111110111","000000000000010000","111111111111101110","111111111111010100","111111111111110101","111111111111101000","111111111111110100","000000000000010110","000000000000001110","000000000000010110","000000000000001100","000000000000001110","000000000000000000","111111111111110010","111111111111111010","000000000000000000","000000000000001111","111111111111110111","111111111111101010","000000000000010010","000000000000000011","111111111111101010","111111111111100111","111111111111101000","000000000000011101","000000000000001110","111111111111110111","000000000000000101"),
("111111111111101111","000000000000010011","111111111111110100","111111111111110110","000000000000000100","000000000000000010","000000000000011110","111111111111101000","000000000000000000","000000000000000101","111111111111110000","111111111111011101","000000000000000001","000000000000000000","000000000000001111","111111111111101100","000000000000001001","111111111111100001","111111111111101011","111111111111100001","000000000000000101","000000000000011111","111111111111101010","000000000000001001","000000000000001110","111111111111101001","000000000000000011","000000000000000111","111111111111111111","111111111111010010","111111111111111000","000000000000001001","000000000000010011","000000000000011010","111111111111101001","111111111111010011","000000000000001100","111111111111110011","111111111111111001","000000000000011100","111111111111110010","000000000000000101","111111111111111001","111111111111110111","000000000000001001","000000000000010001","000000000000001001","000000000000000010","000000000000011000","000000000000001000","000000000000001100","111111111111101100","000000000000001110","000000000000010110","111111111111100111","000000000000001001","000000000000000000","000000000000001011","000000000000011001","111111111111111001","000000000000010010","000000000000000011","111111111111111000","000000000000010110","111111111110100100","000000000000001111","111111111111111010","000000000000000001","000000000000000000","111111111111100111","111111111111110010","111111111111011100","000000000000000010","111111111111111100","111111111111111100","111111111111101010","000000000000010000","000000000000000110","000000000000011000","111111111111110111","111111111111110111","000000000000011110","000000000000010100","000000000000010110","111111111111111101","000000000000000111","000000000000001011","000000000000010100","111111111111110011","000000000000011011","000000000000001011","000000000000001001","111111111111010111","000000000000001001","000000000000001000","111111111111101110","111111111111110011","000000000000100010","000000000000100100","000000000000000110","111111111111111100","000000000000000000","111111111111111110","111111111111110111","111111111111011111","111111111111111001","111111111111111001","000000000000001010","111111111111110111","000000000000011111","111111111111110010","000000000000111000","111111111111101111","111111111111110110","000000000000001101","000000000000000110","111111111111110111","000000000000000010","111111111111111101","000000000000010011","000000000000000000","111111111111111110","111111111111110010","111111111111010110","111111111111111110","000000000000010001","111111111111100001","000000000000000001"),
("111111111111000110","000000000000000100","000000000000000001","111111111111011101","111111111111101111","000000000000001001","000000000000011100","111111111111110110","111111111111110011","000000000000010100","111111111111110111","111111111111110011","111111111111111011","111111111111011101","000000000000011101","111111111111100111","000000000000010101","111111111111011000","111111111111100011","000000000000000011","000000000000001101","000000000000011110","111111111111110010","000000000000011100","000000000000010110","000000000000000110","111111111111111111","111111111111110011","000000000000001101","111111111111010100","111111111111100011","000000000000010111","000000000000000010","000000000000000100","111111111111110111","111111111111100111","111111111111101111","111111111111111100","000000000000000110","000000000000010000","000000000000010110","000000000000011011","000000000000010111","111111111111100111","111111111111111000","000000000000101011","111111111111110010","000000000000001010","111111111111111001","000000000000001101","000000000000010101","111111111111111011","000000000000000000","000000000000011101","000000000000000001","111111111111111010","111111111111011100","000000000000010111","000000000000010100","111111111111110100","000000000000100101","111111111111111011","000000000000000100","000000000000000111","111111111111110011","000000000000001010","111111111111011001","000000000000001101","000000000000011001","111111111111111111","000000000000000011","111111111111110100","111111111111111011","111111111111100101","000000000000000110","111111111111110100","111111111111101010","111111111111111011","000000000000011011","000000000000010000","000000000000001110","111111111111101110","000000000000000010","000000000000100010","111111111111110011","000000000000001011","000000000000001101","000000000000010110","000000000000001000","000000000000100001","000000000000010000","000000000000010010","111111111111111011","000000000000001011","111111111111110011","111111111111010100","000000000000000011","000000000000011010","000000000000001000","111111111111110101","111111111111110101","000000000000011000","000000000000100100","111111111111011001","111111111111100000","111111111111110110","111111111111110110","000000000000010001","111111111111111101","111111111111111111","111111111111100010","000000000000100000","000000000000001101","111111111111110101","111111111111110010","000000000000001001","000000000000001000","000000000000001001","111111111111110011","000000000000011010","000000000000000101","111111111111101111","000000000000001010","111111111111111101","000000000000000011","000000000000011010","111111111111110000","000000000000001001"),
("111111111111000111","000000000000011011","000000000000000110","111111111111011001","000000000000001100","111111111111111110","000000000000011110","111111111111110000","000000000000000101","000000000000001000","111111111111111110","111111111111111000","111111111111011110","111111111111001011","000000000000010010","111111111111111100","000000000000010110","111111111111011101","111111111111100111","000000000000000110","000000000000000110","000000000000000000","111111111111110111","000000000000000010","000000000000001001","111111111111110101","111111111111110010","111111111111111111","000000000000001010","111111111111010111","111111111111101110","000000000000010011","111111111111100100","000000000000000110","111111111111110000","111111111111100100","111111111111111111","111111111111110111","111111111111100101","000000000000000000","000000000000001011","000000000000000111","000000000000001010","111111111111110011","111111111111111001","000000000000101000","000000000000010000","000000000000100010","000000000000000000","111111111111111100","000000000000010010","111111111111110000","111111111111111101","000000000000001110","111111111111111110","111111111111111101","111111111111001100","111111111111111000","000000000000010110","111111111111111011","000000000000001111","000000000000000001","111111111111011100","000000000000000000","111111111111100010","111111111111111111","111111111111100010","111111111111111101","111111111111111101","111111111111110110","111111111111101101","111111111111000010","111111111111011001","111111111111110100","000000000000000101","000000000000011001","000000000000000011","000000000000001111","000000000000001010","000000000000000100","111111111111111011","000000000000000110","000000000000010001","000000000000001100","111111111111011110","111111111111111101","000000000000011100","000000000000001101","111111111111101110","000000000000011001","000000000000001111","000000000000001000","000000000000011111","000000000000010001","000000000000000000","111111111111101001","000000000000010100","000000000000011110","111111111111010010","111111111111100010","000000000000010111","000000000000100000","000000000000000101","111111111111001001","000000000000010010","000000000000011000","111111111111101100","111111111111111110","111111111111100011","000000000000011110","111111111111101111","000000000000110010","111111111111110000","111111111111110001","111111111111110011","000000000000011101","000000000000001001","000000000000000111","111111111111111111","111111111111110111","111111111111110010","000000000000010001","000000000000001101","111111111111110101","000000000000100100","111111111111111011","111111111111110011","111111111111110010"),
("111111111111010101","000000000000110000","111111111111111011","111111111111010010","111111111111110100","111111111111101111","000000000000000000","111111111111111011","111111111111111111","000000000000101100","111111111111101111","000000000000010010","111111111111101010","111111111111101000","000000000000001110","000000000000001010","000000000000010110","111111111111011100","111111111111110011","000000000000001101","000000000000010111","000000000000010011","000000000000000000","000000000000000011","000000000000100111","000000000000000011","000000000000000110","111111111111101001","000000000000011001","000000000000000000","111111111111101111","000000000000010101","111111111111101010","111111111111111111","000000000000000111","111111111111100101","111111111111111111","111111111111110111","111111111111010000","000000000000000101","000000000000011100","111111111111100110","000000000000101101","000000000000000000","111111111111010010","111111111111110101","000000000000110000","000000000000001111","000000000000010011","111111111111110100","000000000000000000","000000000000000001","000000000000000110","000000000000000011","111111111111101111","111111111111100110","111111111111011110","000000000000001010","111111111111111000","111111111111101100","000000000000001010","111111111111111010","111111111111010111","111111111111110110","111111111111111010","000000000000011001","111111111111011111","000000000000011001","000000000000110011","000000000000010101","111111111111101000","111111111111101001","111111111111011000","000000000000010110","111111111111111011","000000000000011101","000000000000000000","111111111111010011","111111111111111010","111111111111111111","111111111111111110","111111111111100100","000000000000000111","111111111111100001","111111111111100111","000000000000000001","000000000000010101","000000000000011000","111111111111100000","000000000000001001","111111111111101101","111111111111110100","000000000000110010","000000000000011000","111111111111110110","111111111111000011","000000000000100010","000000000000000000","111111111110110111","111111111111011111","111111111111110110","000000000000011011","000000000000000010","111111111111011110","000000000000011001","000000000000000011","111111111111011000","000000000000011000","111111111111011101","111111111111111000","111111111111011011","000000000000001011","111111111111111000","111111111111111100","111111111111111000","000000000000000111","000000000000010000","000000000000000010","111111111111101000","000000000000000000","111111111111011100","000000000000001111","000000000000000010","000000000000010010","000000000000100010","000000000000000100","111111111111111100","111111111111101101"),
("111111111111100001","000000000000010111","000000000000001000","111111111111011010","111111111111111101","111111111111111010","111111111111110100","111111111111111110","111111111111111001","000000000001000001","111111111111101110","000000000001000011","111111111111110010","111111111111011000","111111111111010010","000000000000000111","000000000000100010","111111111111011111","000000000000000100","111111111111111110","000000000000010010","000000000000010110","000000000000011001","000000000000000111","000000000000010101","111111111111111000","111111111111100101","111111111111011011","000000000000001111","000000000000010111","000000000000000010","111111111111111000","111111111111100000","000000000000000111","111111111111110101","111111111111110001","000000000000011100","000000000000000111","111111111111101100","000000000000000110","000000000000100001","111111111111110010","000000000000100101","000000000000001110","111111111111100111","111111111111111001","000000000000010101","000000000000000100","000000000000001000","111111111111011101","000000000000011101","000000000000010100","111111111111111101","111111111111111010","111111111111110101","111111111111111001","111111111111010011","111111111111111001","111111111111111110","000000000000000100","111111111111011110","111111111111101010","111111111111011110","111111111111100100","000000000000001000","111111111111110010","111111111111011001","000000000000011101","000000000000101101","000000000000001110","111111111111110100","000000000000000010","111111111111011000","111111111111110110","111111111111110101","000000000000100011","111111111111110100","111111111111011000","111111111111011101","000000000000100001","111111111111101100","111111111111001111","000000000000010000","000000000000000000","000000000000001011","111111111111110011","000000000000010011","000000000000000110","111111111111101100","111111111111110111","000000000000000110","111111111111110110","000000000000100100","000000000000001110","111111111111100100","111111111111011101","000000000000101001","111111111111111010","111111111111101001","111111111110111000","000000000000011001","000000000000010011","111111111111001101","111111111111101110","111111111111110101","000000000000010011","111111111111110101","000000000000000010","111111111111011001","111111111111111101","111111111111001011","000000000000001110","111111111111111111","000000000000000101","111111111111110101","000000000000010100","000000000000010011","111111111111111001","111111111111110010","000000000000000111","111111111111110011","000000000000110000","000000000000010000","111111111111001110","000000000000011100","111111111111101010","000000000000000001","111111111111111100"),
("111111111111110100","000000000000000011","000000000000000000","000000000000001100","111111111111110011","000000000000001001","000000000000101010","000000000000011001","000000000000010111","000000000000001100","000000000000010000","000000000000001100","111111111111001111","111111111111010011","111111111111100011","000000000000101001","000000000000010011","000000000000000101","111111111111111100","000000000000000011","000000000000000101","111111111111111100","000000000000001101","111111111111111110","111111111111011100","000000000000000011","111111111111110100","111111111111110100","111111111111110110","000000000000010000","111111111111101101","111111111111111010","111111111111110010","111111111111101001","111111111111100101","000000000000001111","111111111111110101","000000000000000110","111111111111101011","111111111111110101","111111111111111000","111111111111110110","000000000000001111","000000000000010111","111111111111111011","111111111111110011","000000000000000110","000000000000000110","111111111111010110","111111111111111010","000000000000100100","000000000000010000","111111111111110101","111111111111011101","000000000000011111","000000000000001110","111111111111110100","111111111111101111","111111111111101001","111111111111111111","111111111111100010","000000000000001001","000000000000001100","000000000000001000","111111111111101010","111111111111010110","111111111111011000","000000000000000011","000000000000011010","111111111111011010","000000000000011001","000000000000000000","111111111111000010","000000000000011011","000000000000010001","000000000000010101","000000000000000101","111111111111011000","111111111111101111","000000000000110111","111111111111101100","111111111111110110","000000000000110111","111111111111111101","111111111111011110","111111111111100000","111111111111110101","000000000000000001","111111111111001110","111111111111111011","111111111111101111","111111111111110100","111111111111111110","000000000000001000","000000000000010001","111111111111101100","000000000000110011","111111111111100110","111111111111011001","111111111111110010","000000000000101111","000000000000000111","111111111111010001","111111111111111011","000000000000001001","000000000000011111","000000000000001110","111111111111110101","000000000000001010","111111111111110011","111111111111110001","111111111111111111","111111111111111010","000000000000001001","111111111111110101","111111111111110101","111111111111111001","111111111111100101","111111111111100101","111111111111101100","111111111111100010","000000000000110001","000000000000010110","000000000000100010","000000000000100000","000000000000001101","111111111111110101","000000000000001011"),
("000000000000101011","111111111111110000","111111111111100000","000000000000010100","111111111111101000","000000000000011110","000000000000100100","111111111111111110","000000000000010100","111111111111110101","000000000000100001","111111111111001010","000000000000001111","111111111111111110","111111111111110111","000000000000001110","000000000000001011","000000000000001101","111111111111110000","000000000000001001","000000000000110100","000000000000001000","000000000000011010","111111111111010111","111111111111100100","000000000000111100","111111111111001011","000000000000000110","111111111111110000","111111111111100111","000000000000101111","111111111111100101","000000000000011110","111111111111101010","000000000001010001","111111111111110000","000000000000011001","000000000000011111","111111111111101110","000000000000000101","111111111111111000","111111111111011001","000000000000110110","000000000000111011","111111111111011101","111111111111100000","000000000000011111","000000000000111010","111111111111001101","111111111111101000","000000000000000101","000000000000011101","111111111111001110","000000000000101101","000000000000011011","000000000000101111","111111111111011110","000000000000011110","111111111111000110","000000000000001101","111111111111101010","000000000000010101","000000000000010011","111111111111110110","111111111111011010","111111111111100000","111111111111010000","111111111111111001","000000000000101100","000000000000000000","000000000000011001","111111111111110100","111111111111011111","000000000000100011","111111111111101101","000000000000101110","000000000000111111","000000000000001010","111111111111101001","000000000000110100","111111111111100001","000000000000011101","000000000000110110","111111111111110101","000000000000010001","111111111111100101","000000000000001101","000000000000001011","111111111111010011","111111111111101010","111111111111011011","111111111111100100","111111111111010011","000000000000101000","111111111111100111","111111111111110011","111111111111101111","000000000000010111","111111111111100101","111111111111101000","000000000000110001","111111111111101010","111111111111101110","000000000000011100","111111111111111111","000000000000011000","111111111111100101","111111111111010010","111111111111000100","111111111111010101","111111111111111101","000000000000001101","111111111111100101","111111111111100001","000000000000010010","000000000000111111","000000000000001000","000000000000011000","111111111111010010","000000000000000000","000000000000100000","000000000000110011","000000000000101110","000000000000000100","000000000000010110","111111111111110000","000000000000101111","111111111111110010"),
("000000000000010101","111111111111100111","000000000000000100","111111111111111111","111111111111111001","000000000000011001","000000000000011010","000000000000010010","000000000000010111","000000000000001010","000000000000001100","111111111111100101","000000000000000111","000000000000000000","111111111111101100","111111111111111000","000000000000000011","000000000000011011","111111111111111001","000000000000011100","000000000000010001","111111111111101101","000000000000000000","111111111111101001","111111111111100011","000000000000010101","111111111111111100","111111111111111111","111111111111111101","000000000000001001","111111111111111110","111111111111110011","111111111111111011","111111111111111101","000000000000011101","111111111111111111","111111111111111100","000000000000001110","000000000000000111","000000000000001010","111111111111101000","111111111111110010","000000000000011110","000000000000000100","111111111111100000","000000000000001010","000000000000000010","111111111111111101","111111111111100101","111111111111110110","000000000000000111","000000000000000011","000000000000000110","000000000000011001","000000000000000010","000000000000001000","111111111111101010","111111111111101101","000000000000000011","000000000000000011","111111111111110010","000000000000010000","111111111111110100","000000000000000000","000000000000010000","111111111111100010","000000000000001110","111111111111110001","000000000000011000","000000000000000110","000000000000000101","111111111111111101","111111111111110001","000000000000000100","111111111111110101","111111111111111111","000000000000011000","000000000000010000","111111111111100100","000000000000011111","000000000000000101","000000000000001000","000000000000010010","111111111111100100","000000000000001001","000000000000000011","111111111111110110","000000000000001011","111111111111101110","111111111111110101","000000000000000001","000000000000001001","000000000000000111","000000000000100011","000000000000010011","111111111111111101","111111111111110100","000000000000010001","111111111111100101","111111111111110000","000000000000000010","111111111111100011","111111111111111110","000000000000001001","111111111111110100","000000000000000110","000000000000000101","000000000000000000","000000000000000101","111111111111101011","111111111111110111","111111111111111001","111111111111101011","111111111111110101","000000000000000111","000000000000011010","111111111111111101","111111111111111101","000000000000000001","111111111111110001","000000000000010101","111111111111111010","000000000000000000","111111111111111101","000000000000010111","000000000000001011","000000000000001101","000000000000001000"),
("000000000000000111","111111111111110001","000000000000001110","000000000000000000","000000000000001000","111111111111101101","111111111111101010","000000000000000010","111111111111110111","111111111111101111","000000000000001001","000000000000000111","111111111111111011","000000000000001111","111111111111100101","111111111111110110","000000000000001101","000000000000001100","111111111111111101","111111111111111100","000000000000000100","111111111111110111","000000000000001000","000000000000000000","000000000000000000","111111111111111110","111111111111101101","000000000000000011","111111111111111011","000000000000000011","000000000000000100","111111111111111000","111111111111111000","000000000000010010","111111111111110010","000000000000001101","111111111111110111","000000000000001010","111111111111101110","000000000000010110","000000000000001010","111111111111111011","111111111111111001","111111111111101010","111111111111101101","111111111111110011","111111111111111110","111111111111110110","000000000000010110","111111111111101101","111111111111111000","000000000000001011","000000000000000111","000000000000010011","000000000000000000","000000000000001011","111111111111111111","111111111111111100","000000000000001100","111111111111111101","000000000000000100","111111111111111111","111111111111110011","111111111111101000","111111111111100111","000000000000010010","000000000000001001","000000000000000000","111111111111111001","000000000000000111","111111111111110000","111111111111111000","111111111111110010","000000000000001001","111111111111110100","111111111111101110","000000000000000101","111111111111110101","000000000000000111","111111111111111001","000000000000010000","000000000000000000","000000000000001100","111111111111110001","111111111111111010","000000000000001000","000000000000000000","000000000000010010","111111111111111001","000000000000000101","000000000000001100","111111111111101011","111111111111101011","000000000000001110","000000000000001001","111111111111110110","000000000000000100","111111111111111001","000000000000010110","111111111111111111","000000000000001111","000000000000001111","111111111111101000","000000000000001001","111111111111110101","000000000000010001","000000000000000010","000000000000000001","000000000000001010","000000000000001101","000000000000000001","000000000000001110","000000000000001001","111111111111111011","000000000000000010","111111111111100111","000000000000001010","111111111111110011","111111111111111100","000000000000000000","000000000000000000","111111111111111100","000000000000001111","000000000000001010","111111111111110100","111111111111111010","111111111111111110","111111111111101111"),
("111111111111110101","111111111111111000","111111111111111010","000000000000000110","000000000000000101","000000000000000010","111111111111110000","111111111111111010","000000000000001110","000000000000000110","000000000000000100","000000000000000000","000000000000000110","111111111111111111","000000000000001011","000000000000000001","000000000000100101","000000000000000100","000000000000001011","000000000000010101","000000000000010000","000000000000000010","000000000000010110","000000000000000011","111111111111110010","111111111111110101","111111111111111101","111111111111101100","000000000000010101","000000000000001000","000000000000000100","000000000000010100","000000000000011001","000000000000001010","111111111111111111","000000000000011000","111111111111101111","000000000000001001","000000000000010100","000000000000000111","000000000000010000","111111111111100101","111111111111111101","111111111111111101","000000000000001111","000000000000000011","111111111111110001","000000000000000000","000000000000011011","000000000000000110","111111111111110000","000000000000001100","111111111111111100","111111111111111100","000000000000000000","000000000000000100","000000000000010001","000000000000011000","000000000000000000","000000000000010011","000000000000000101","111111111111101010","000000000000001001","111111111111111000","111111111111110000","111111111111111001","000000000000000010","111111111111111011","000000000000000110","111111111111101011","000000000000000110","000000000000011010","111111111111110000","000000000000010011","111111111111111000","000000000000000111","111111111111110010","000000000000000100","111111111111110010","111111111111111001","000000000000010100","000000000000000010","111111111111100110","000000000000011101","111111111111111010","000000000000000010","111111111111111110","000000000000000000","000000000000000010","000000000000000000","111111111111101011","000000000000011010","111111111111111010","000000000000001010","111111111111111111","111111111111111001","111111111111111010","000000000000001111","000000000000011101","000000000000000010","111111111111101111","000000000000000000","000000000000010100","111111111111111000","000000000000001010","000000000000001011","000000000000011011","000000000000001111","000000000000100000","111111111111110101","111111111111110001","111111111111110100","111111111111111110","000000000000000000","000000000000011001","000000000000000101","000000000000001000","111111111111110101","000000000000001000","000000000000010011","111111111111100100","111111111111101010","000000000000001010","111111111111110101","000000000000000000","111111111111110110","111111111111110011","000000000000010001"),
("000000000000010101","000000000000010010","000000000000000011","000000000000001011","000000000000011010","000000000000010100","111111111111000110","000000000000100001","111111111111111001","000000000000011111","000000000000001100","000000000000010100","000000000000000101","111111111111111111","111111111111101110","111111111111101101","000000000000100100","000000000000000001","000000000000010000","000000000000001100","000000000000000101","000000000000010011","000000000000110111","000000000000010000","111111111111101010","111111111111110010","000000000000101000","111111111111010001","000000000000010100","000000000000011001","111111111111111001","000000000000001111","111111111111101000","111111111111110101","111111111111111000","000000000000100001","111111111111100101","000000000000110011","000000000000000110","000000000000101001","111111111111111001","000000000000000101","000000000000000110","000000000000100001","000000000000000100","000000000000000111","111111111111111100","000000000000010111","000000000000000100","000000000000000101","000000000000000001","000000000000010111","111111111111111001","111111111111010010","111111111111111111","111111111111101110","111111111111111110","000000000000001010","111111111111011010","000000000000001100","000000000000000110","000000000000000010","111111111111011000","000000000000011010","000000000000011001","111111111111010001","111111111111100101","000000000000010101","111111111111101011","000000000000100010","111111111111110111","000000000000010111","111111111111101101","111111111111100101","000000000000011101","111111111111111100","111111111111101010","111111111111110100","111111111111111100","111111111111110011","000000000000010101","111111111111110010","000000000000011110","000000000000001001","000000000000011001","000000000000000011","000000000000011001","000000000000110011","000000000000001101","111111111111110000","000000000000100010","111111111111111010","111111111111011111","111111111111111110","111111111111011101","111111111111111101","000000000000001100","111111111111011101","111111111111111010","000000000000001011","000000000000000100","000000000000100101","111111111111101001","000000000000001100","111111111111110001","000000000000001110","111111111111011111","111111111111011001","000000000000001000","111111111111111100","111111111111011011","111111111111010000","000000000000110011","000000000000010111","000000000000000100","111111111111101011","111111111111100010","000000000000001111","111111111111111011","000000000000011111","000000000000010101","000000000000001110","111111111111110111","000000000000110111","000000000000000100","111111111111001111","111111111111110111","000000000000000000"),
("111111111111101111","111111111111101101","000000000000010001","000000000000010010","000000000000000101","000000000000101001","000000000000001010","111111111111111011","000000000000000110","000000000000000010","111111111111101000","111111111111100001","111111111111111100","111111111111110110","000000000000100011","111111111111111111","000000000000100111","000000000000000010","000000000000011010","000000000000000100","111111111111111011","000000000000001000","111111111111101000","000000000000000000","111111111111011011","000000000000010001","000000000000001100","000000000000001111","000000000000000111","111111111111110000","000000000000001110","111111111111111010","111111111111110100","111111111111010100","000000000000010011","111111111111111111","111111111111111101","111111111111111000","000000000000000000","000000000000001110","111111111111011111","000000000000010000","000000000000101011","111111111111111011","000000000000000001","111111111111111110","111111111111101101","000000000000101000","111111111111101011","111111111111101110","000000000000000000","000000000000010100","111111111111110011","111111111111100100","000000000000101011","000000000001001100","111111111111100100","111111111111111110","111111111111111000","111111111111110001","111111111111100000","000000000000101001","000000000000011110","000000000000000101","111111111111110001","111111111111111100","111111111111110100","111111111111010100","111111111111011000","000000000000001010","111111111111110100","111111111111101010","111111111111110011","000000000000010110","000000000000000000","111111111111111000","000000000000011010","111111111111110100","000000000000100101","000000000000010001","111111111111101101","111111111111110000","000000000000101110","111111111111101011","111111111111111010","111111111111110001","000000000000111001","000000000000001111","000000000000000000","000000000000100011","111111111111111110","111111111111100000","000000000000001000","111111111111100011","111111111111111101","111111111111101111","000000000000001000","000000000000011111","111111111111100011","000000000000000110","000000000000010001","111111111111111010","111111111111010100","111111111111010010","111111111111110111","111111111111111000","000000000000011011","111111111111100000","111111111111110111","111111111111101001","111111111111111010","000000000000010111","111111111111110101","000000000000001011","000000000000110111","111111111111101101","111111111111110111","111111111111110001","111111111111101101","000000000000000100","111111111111100010","000000000000010000","000000000000001011","000000000000011111","000000000000010000","111111111111001001","111111111111101001","111111111111101111"),
("000000000000010011","000000000000001001","000000000000000111","000000000000001101","000000000000110100","000000000000000101","111111111111011111","000000000000010110","111111111111100001","000000000000000101","111111111111000010","000000000000000111","111111111111001011","000000000000000010","000000000000001001","111111111111100111","000000000000001000","000000000000000010","111111111111111000","111111111111110110","111111111111111000","111111111111101110","000000000000001000","111111111111101100","000000000000011000","111111111111110110","111111111111111011","000000000000010011","000000000000000100","111111111111110010","111111111111111011","111111111111011010","000000000000100010","111111111111010010","111111111111100110","111111111111000001","111111111111111011","111111111111111001","111111111111011000","000000000000010110","000000000000010001","111111111111111101","111111111111110100","111111111111100101","000000000000001101","111111111111101101","111111111111010001","000000000000010100","111111111111111100","000000000000000010","111111111111100001","000000000000100000","111111111111111110","111111111111011011","111111111111111010","000000000000100000","111111111111110010","000000000000000001","000000000000000000","111111111111111010","111111111111111100","000000000000111100","000000000000010001","111111111111111110","000000000000001100","000000000000001010","111111111111111011","111111111111101011","111111111111011101","111111111111110100","111111111111100011","111111111111110101","000000000000001101","000000000000000111","111111111111011010","111111111111010110","111111111111111110","000000000000001010","111111111111111000","111111111111100101","111111111111111001","000000000000100000","000000000000011011","000000000000011011","111111111111111010","000000000000000000","000000000000001011","000000000000000101","111111111111101010","000000000000010110","000000000000000010","000000000000001111","000000000000000001","000000000000001010","000000000000001110","111111111111101011","000000000000000000","000000000000001100","000000000000010100","111111111111111110","000000000000010010","111111111111111101","000000000000010110","111111111111010110","111111111111100111","111111111111111000","111111111111101111","111111111111001101","000000000000000000","000000000000000010","111111111111110111","000000000000011100","111111111111110000","111111111111111010","000000000000010010","000000000000010001","111111111111101101","000000000000010001","111111111111011101","000000000000000100","111111111111101001","000000000000000110","000000000000001111","111111111111111001","000000000000001100","111111111111010101","111111111111101111","000000000000000010"),
("000000000000100010","000000000000101011","000000000000010111","000000000000001010","000000000000001101","000000000000010101","111111111111101111","111111111111111100","111111111111001100","000000000000010001","111111111111000010","111111111111110000","111111111111001000","000000000000000111","000000000000001010","111111111111101100","000000000000010001","111111111111100010","111111111111010110","111111111111110100","000000000000010000","111111111111111111","000000000000001110","111111111111101011","000000000000001111","111111111111111000","000000000000010101","000000000000001010","000000000000010100","111111111111100000","111111111111110101","111111111111101000","111111111111110110","111111111111110100","111111111111110001","111111111111001011","111111111111101110","111111111111101000","111111111111101000","000000000000100010","000000000000000101","111111111111110010","111111111111101100","111111111111010000","000000000000001111","111111111111101010","111111111111101111","000000000000001010","111111111111101110","111111111111111100","000000000000011110","000000000000100000","000000000000000000","111111111111100000","111111111111010111","000000000000001100","111111111111011101","000000000000011101","000000000000010010","000000000000010000","000000000000100011","000000000001010100","111111111111111100","111111111111111110","111111111111110011","000000000000001011","000000000000001000","111111111111111011","111111111111100110","000000000000001101","000000000000000001","111111111111101101","000000000000110000","111111111111111010","111111111111011100","111111111111110001","000000000000000111","111111111111110011","111111111111101001","000000000000010001","111111111111111100","000000000000000101","000000000000000101","111111111111100010","111111111111110110","111111111111101011","111111111111111111","111111111111111000","111111111111101111","000000000000000110","111111111111110011","111111111111110111","000000000000010010","000000000000010111","111111111111110101","111111111111110101","111111111111111011","000000000000000010","000000000000000000","111111111111110110","000000000000010010","000000000000000011","000000000000000001","111111111111100100","111111111111101010","000000000000100011","111111111111111110","111111111111111111","111111111111010111","111111111111110101","111111111111011010","000000000000010010","000000000000001101","111111111111101000","111111111111110011","000000000000110010","000000000000001011","000000000000000000","111111111111100011","111111111111011000","111111111111010110","111111111111011111","111111111111111010","111111111111110011","000000000000001100","111111111111111100","111111111111101010","111111111111110111"),
("000000000000001111","000000000000101110","000000000000100111","000000000000010100","111111111111110011","000000000000010000","000000000000001111","000000000000000000","111111111111010100","000000000000110010","111111111110110000","111111111111110010","111111111111011111","111111111111111010","000000000000001110","000000000000010011","000000000000101100","000000000000000111","111111111111100010","111111111111101010","000000000000010000","000000000000000010","111111111111111100","111111111111100101","111111111111110110","111111111111111100","000000000000000011","111111111111101100","111111111111111100","111111111111110101","000000000000011000","000000000000000010","111111111111101010","111111111111010110","111111111111101001","111111111111101100","000000000000001111","111111111111111101","111111111111100010","000000000000001100","111111111111100010","000000000000000010","111111111111100000","111111111111001001","000000000000011110","000000000000000101","111111111111110011","000000000000010111","000000000000001110","111111111111011101","000000000000001000","000000000000011111","111111111111111001","111111111111101101","111111111111000001","000000000000010100","111111111111010110","000000000000000000","000000000000010001","000000000000000011","111111111111111000","000000000001001000","000000000000000000","111111111111111000","111111111111011110","000000000000001000","000000000000100100","000000000000000110","111111111111001111","000000000000000100","000000000000010111","111111111111110000","000000000000110001","000000000000000000","000000000000001011","111111111111110010","111111111111111101","000000000000001101","000000000000001101","111111111111111011","111111111111110001","000000000000000000","000000000000001100","111111111111101111","111111111111111010","111111111111111011","000000000000010000","111111111111110111","111111111111100110","111111111111111101","000000000000000100","111111111111101011","111111111111110011","111111111111111110","111111111111111000","111111111111101101","000000000000001100","000000000000001100","111111111111011100","111111111111111001","000000000000001010","111111111111110001","000000000000000001","111111111111101101","111111111111100001","000000000000001101","111111111111110001","000000000000000000","111111111111010100","000000000000000111","111111111111111011","000000000000001111","000000000000001101","111111111111111010","000000000000000000","000000000000011011","111111111111111101","111111111111001110","111111111111001101","111111111111000110","111111111111001001","111111111111111010","111111111111101111","111111111111110101","111111111111111010","111111111111101100","111111111111011001","111111111111110111"),
("000000000000100100","000000000000111101","000000000000011111","000000000000000001","000000000000001101","000000000000010001","000000000000000010","000000000000011100","111111111111100000","000000000000100011","111111111110111001","000000000000001010","111111111111100000","000000000000010010","000000000000010010","000000000000000000","000000000000001011","111111111111111100","111111111111011101","000000000000000101","111111111111101100","000000000000100100","000000000000011101","111111111111110101","111111111111111111","111111111111111111","000000000000001001","000000000000001101","111111111111111100","111111111111011011","111111111111110001","111111111111101001","111111111111100111","111111111111101111","111111111111100011","111111111111011111","000000000000000100","111111111111101010","111111111111100001","000000000000000010","111111111111110101","111111111111110100","111111111111110111","111111111111100110","000000000000010101","111111111111111111","111111111111111111","000000000000101100","000000000000001001","000000000000000101","000000000000000111","000000000000001110","000000000000010000","111111111111010011","111111111111010011","000000000000001000","111111111111001011","000000000000000101","000000000000000110","000000000000000111","111111111111111101","000000000000010000","000000000000001111","000000000000010000","111111111110100110","000000000000001101","000000000000011101","111111111111111011","000000000000010000","000000000000010001","111111111111101101","111111111111110110","000000000000100010","111111111111101101","111111111111110111","111111111111101010","111111111111110100","111111111111101111","000000000000011011","000000000000011111","000000000000011001","111111111111111010","000000000000010110","111111111111110000","111111111111110110","000000000000001000","111111111111111100","111111111111101011","000000000000010101","000000000000000011","000000000000011101","000000000000000110","000000000000000011","000000000000100001","000000000000000010","111111111111101011","000000000000000001","111111111111110100","111111111111101101","000000000000000101","000000000000010011","000000000000000100","111111111111111111","111111111111101101","111111111111111010","000000000000000110","000000000000100000","111111111111110011","000000000000000010","000000000000000101","111111111111110011","111111111111100111","000000000000001011","111111111111111110","000000000000001111","000000000000001100","000000000000001000","111111111111000000","111111111111011100","111111111111100100","111111111111100100","111111111111011110","111111111111110011","000000000000000011","000000000000010100","111111111111110100","111111111111110111","111111111111101100"),
("000000000000100100","000000000000101010","000000000000100101","000000000000001100","000000000000001001","000000000000010011","000000000000010101","000000000000010110","111111111111011011","000000000000011000","111111111110100000","000000000000001011","111111111111111010","000000000000110001","111111111111111110","000000000000011001","111111111111111110","000000000000000010","111111111111001010","111111111111110011","111111111111110111","000000000000010110","000000000000011001","111111111111101111","111111111111111111","000000000000000111","111111111111111011","111111111111111010","000000000000001101","111111111111111101","111111111111111000","000000000000000001","111111111111110010","000000000000000000","111111111111111010","111111111111100101","111111111111101101","111111111111101101","111111111111110101","111111111111110111","111111111111001101","000000000000000010","111111111111011010","000000000000001001","000000000000010000","000000000000011001","111111111111001000","000000000000110110","111111111111110000","000000000000010010","000000000000100011","000000000000001100","111111111111101100","111111111111110011","111111111111001001","000000000000100001","111111111111100110","000000000000000001","000000000000011110","111111111111111100","111111111111110110","000000000000001000","000000000000100111","000000000000011100","111111111111010101","000000000000001010","111111111111111001","111111111111110101","000000000000110000","000000000000010001","111111111111111111","111111111111111000","000000000000000011","000000000000001101","111111111111111111","111111111111100010","111111111111111101","000000000000000010","000000000000010001","000000000000011010","000000000000001001","111111111111111011","000000000000100000","111111111111110000","000000000000000101","000000000000010110","111111111111111001","111111111111110100","000000000000000100","000000000000011111","000000000000000101","000000000000000001","000000000000001101","000000000000100101","111111111111111011","111111111111111111","111111111111111110","000000000000000100","111111111111101101","000000000000001001","000000000000100001","000000000000001001","111111111111111101","111111111111111010","111111111111101000","000000000000011111","000000000000100001","111111111111100111","000000000000001001","000000000000001101","000000000000001101","111111111111111011","000000000000011111","111111111111111000","000000000000011000","111111111111111101","000000000000000110","111111111111000101","000000000000000011","111111111111101011","111111111111100111","000000000000000001","111111111111101000","111111111111111011","000000000000000010","000000000000001001","111111111111101111","111111111111101111"),
("111111111111111001","111111111111110111","000000000000111111","111111111111111111","000000000000100010","000000000000001111","000000000000001101","000000000000011101","111111111111110101","111111111111110010","111111111110010110","000000000000011010","111111111111011001","000000000000000111","111111111111111011","000000000000000001","000000000000010011","000000000000000010","111111111111001011","000000000000000110","000000000000010010","111111111111111111","111111111111111010","111111111111101111","000000000000001000","111111111111110011","111111111111111001","111111111111110011","000000000000000111","111111111111111001","111111111111101110","111111111111110000","111111111111011110","111111111111111100","000000000000000100","111111111111101011","111111111111110100","111111111111100101","000000000000000110","111111111111011000","111111111111100101","111111111111101111","111111111111110101","111111111111111111","000000000000000110","000000000000010010","111111111110111011","000000000000011101","000000000000001001","000000000000000011","000000000000111010","000000000000000000","000000000000011011","111111111111111011","111111111111011101","111111111111111111","000000000000000100","111111111111110101","000000000000000110","000000000000001101","111111111111100110","000000000000001011","000000000000100000","000000000000000010","111111111111111011","000000000000001101","111111111111100011","000000000000000110","000000000000100001","000000000000100000","000000000000001100","000000000000000110","111111111111100100","111111111111110100","111111111111100100","000000000000000010","000000000000010100","111111111111110100","000000000000000110","111111111111111000","111111111111111111","111111111111111000","000000000000100100","111111111111111011","111111111111101100","000000000000010110","000000000000011100","111111111111111011","000000000000011111","000000000000001101","000000000000101100","111111111111110000","000000000000010010","000000000000000000","111111111111111011","111111111111100110","111111111111101000","111111111111100110","111111111111110011","111111111111110010","000000000000010110","111111111111111000","000000000000000011","111111111111111001","111111111111101011","000000000000001001","000000000000100001","111111111111101000","111111111111111010","111111111111111101","111111111111101110","111111111111101111","000000000000000010","111111111111010001","000000000000011011","000000000000001011","111111111111110010","111111111111100000","111111111111110110","111111111111111111","111111111111101110","000000000000010001","111111111111101101","111111111111101011","000000000000100001","111111111111111110","000000000000001000","111111111111111001"),
("000000000000001010","111111111111110111","000000000000100110","111111111111101000","111111111111111000","000000000000000000","000000000000010010","111111111111110111","111111111111011000","000000000000001010","111111111110111100","000000000000010101","111111111111101100","000000000000010001","000000000000000111","000000000000011100","000000000000101001","000000000000000100","111111111111001110","000000000000001001","000000000000000000","111111111111010011","111111111111101010","111111111111111111","000000000000011001","000000000000000110","000000000000010010","111111111111100111","111111111111101000","000000000000011111","111111111111100011","000000000000000001","111111111111111011","111111111111111010","111111111111110001","111111111111110101","000000000000000111","111111111111001101","000000000000110101","111111111111111000","111111111111011100","111111111111111100","000000000000001001","000000000000010110","000000000000000010","000000000000000111","111111111111011101","000000000000011101","000000000000001010","000000000000000100","000000000000110010","111111111111110100","000000000000010000","000000000000000111","111111111111011011","000000000000001100","000000000000000100","111111111111101001","000000000000000110","000000000000001001","111111111111101000","000000000000010100","000000000000100001","000000000000010001","000000000000010110","000000000000100000","000000000000000000","000000000000001000","000000000001001001","000000000000001010","111111111111101000","111111111111101000","111111111111110001","111111111111101100","111111111111100111","000000000000001000","000000000000000010","111111111111100010","000000000000011110","111111111111111101","000000000000000000","000000000000001101","111111111111111101","000000000000000010","111111111111101001","000000000000010001","000000000000011100","000000000000000000","000000000000011111","000000000000001011","000000000000010010","111111111111111100","000000000000001011","111111111111111101","111111111111101110","000000000000010010","111111111111000101","000000000000000010","111111111111100101","111111111111100010","000000000000100110","000000000000010111","111111111111110001","111111111111110011","111111111111111011","000000000000010001","000000000000010001","111111111111111011","000000000000001101","000000000000100101","111111111111110101","111111111111100000","111111111111111011","111111111111111100","000000000000011100","000000000000000100","000000000000000100","111111111111101101","000000000000011100","111111111111110001","111111111111110011","000000000000010100","111111111111100101","111111111110111100","000000000000011111","000000000000001010","000000000000001010","111111111111101110"),
("000000000000000111","111111111111001011","000000000000100001","111111111111111101","000000000000001010","000000000000011000","000000000000001001","111111111111100000","000000000000001100","111111111111001001","111111111111110011","000000000000101111","111111111111101100","111111111111111101","000000000000000101","000000000000010101","000000000000011111","000000000000001010","111111111111011010","111111111111111111","111111111111110011","111111111111011101","111111111111100000","111111111111011111","000000000000001010","000000000000001010","000000000000000000","111111111111110110","111111111111110110","000000000000000000","111111111111110111","000000000000000011","000000000000000111","111111111111101110","111111111111110000","111111111111110010","111111111111111111","111111111111011101","000000000000011111","000000000000000011","111111111111110111","111111111111111001","000000000000101011","000000000000010010","000000000000011010","111111111111110001","000000000000101100","111111111111110110","111111111111111100","111111111111110100","000000000000010011","000000000000000110","000000000000010000","111111111111101101","111111111111100100","111111111111111011","000000000000000110","111111111111101000","111111111111110101","111111111111110000","000000000000000110","111111111111111111","000000000000000110","000000000000011101","000000000000001011","000000000000001100","111111111111110001","111111111111111111","000000000000111010","111111111111101001","000000000000000011","111111111111100111","111111111111110110","000000000000000010","111111111111110010","000000000000011101","000000000000011001","000000000000000000","111111111111111000","000000000000010100","111111111111111011","000000000000000000","000000000000001001","000000000000011001","111111111111110010","000000000000100001","000000000000010000","111111111111110010","000000000000000000","000000000000010010","000000000000011001","000000000000000110","000000000000010000","000000000000011111","111111111111110000","111111111111111110","111111111111001001","000000000000011101","111111111111111111","000000000000000101","000000000000100010","000000000000001000","111111111111110000","000000000000000001","000000000000000010","000000000000011110","000000000000011011","000000000000000000","000000000000011100","000000000000011111","111111111111111010","111111111111101101","000000000000011001","111111111111110001","000000000000100011","000000000000001100","000000000000011101","111111111111110100","000000000000011101","111111111111101100","111111111111100010","000000000000101010","111111111111110010","111111111110001000","000000000000100111","000000000000000011","000000000000100011","111111111111110000"),
("000000000000000000","111111111111000111","000000000000100000","000000000000010111","000000000000000001","000000000000010100","000000000000001010","111111111111011100","111111111111110010","111111111111100011","000000000000011011","000000000000100000","111111111111110110","111111111111110000","111111111111100011","000000000000010010","000000000000001111","111111111111111100","111111111111110010","111111111111110100","000000000000001101","111111111111110111","111111111111101000","111111111111110001","111111111111110011","111111111111111111","000000000000010100","111111111111101010","000000000000000000","000000000000011000","111111111111111110","111111111111101000","111111111111111010","000000000000001010","000000000000000100","000000000000011010","000000000000000110","111111111111111110","000000000000100001","111111111111110000","111111111111100111","000000000000010000","000000000000010100","000000000000001101","000000000000010101","111111111111110010","000000000001000000","111111111111111011","000000000000001001","000000000000001001","111111111111110101","000000000000001101","000000000000001000","000000000000000110","111111111111110011","111111111111110100","000000000000000110","111111111111101001","111111111111101001","111111111111110100","111111111111110001","000000000000000000","111111111111101101","000000000000100010","000000000000110011","000000000000000010","000000000000001110","000000000000101001","000000000000101110","111111111111010011","000000000000010110","111111111111111010","000000000000011011","111111111111101001","111111111111011011","000000000000011010","111111111111111010","111111111111101000","111111111111101111","000000000000000110","000000000000011001","000000000000011010","000000000000001100","000000000000011000","000000000000000001","000000000000010010","000000000000000100","000000000000001100","000000000000000011","111111111111111101","111111111111101001","000000000000000001","000000000000000000","111111111111110010","111111111111111110","000000000000000010","111111111111011101","111111111111110010","000000000000100000","000000000000010010","000000000000101001","111111111111111111","000000000000001011","000000000000100000","000000000000000100","000000000000100101","000000000000000010","111111111111111010","000000000000001101","111111111111110101","111111111111110110","111111111111010100","000000000000101110","000000000000010111","000000000000011101","000000000000100010","000000000000000001","111111111111111101","000000000000101111","111111111111101110","111111111111101000","000000000000001001","111111111111111011","111111111101101001","000000000000101011","111111111111110010","000000000000001011","111111111111110101"),
("000000000000001001","111111111111100111","111111111111110001","000000000000000011","111111111111111101","000000000000011001","111111111111111010","111111111111111000","000000000000100010","111111111110111101","000000000000011011","111111111111111010","000000000000000001","000000000000001110","111111111111101000","000000000000001101","000000000000011101","000000000000001010","111111111111111100","000000000000000010","000000000000000000","000000000000000010","111111111111101000","000000000000101001","111111111111100011","000000000000011101","000000000000001001","000000000000010001","000000000000001001","111111111111101101","000000000000000001","000000000000000011","111111111111110000","111111111111111111","000000000000010011","000000000000001101","111111111111110000","000000000000000100","000000000000011111","000000000000001000","111111111111100001","000000000000010001","000000000000011011","000000000000011001","000000000000011110","111111111111100101","000000000001010010","000000000000010101","000000000000000000","000000000000001010","111111111111001110","111111111111111101","111111111111100100","000000000000001011","111111111111110101","111111111111111111","111111111111110010","111111111111100111","111111111111111000","000000000000000111","111111111111111001","111111111111110010","111111111111110011","000000000000011000","000000000000010011","111111111111011011","111111111111110110","000000000000100010","000000000000100111","111111111111100000","000000000000101110","000000000000010110","111111111111110110","111111111111110010","000000000000001101","111111111111101111","000000000000001110","000000000000010010","111111111111110001","000000000000000010","111111111111110111","000000000000001001","000000000000010100","000000000000110000","000000000000001100","111111111111011001","000000000000001011","111111111111111000","111111111111111010","000000000000011000","111111111111110001","000000000000010100","000000000000001100","111111111111111010","111111111111110100","000000000000000100","111111111111100001","000000000000001010","000000000000001111","000000000000001000","000000000000110010","000000000000010110","000000000000000101","000000000000011000","000000000000100110","000000000000000111","000000000000010000","000000000000010000","000000000000011001","111111111111010111","000000000000000101","000000000000000000","000000000000100100","000000000000000000","000000000000110100","000000000000000110","000000000000000101","111111111111110001","000000000000011000","111111111111111010","111111111111110000","000000000000000010","000000000000011100","111111111110011100","000000000000010101","000000000000000000","000000000000000111","111111111111111001"),
("000000000000101000","111111111111111010","111111111111101011","000000000000001110","000000000000000101","000000000000100010","000000000000001110","000000000000000010","000000000000110010","111111111111110110","000000000000100110","000000000000010100","111111111111111101","000000000000001001","111111111111011010","000000000000001101","111111111111110010","000000000000010001","000000000000010101","111111111111110000","000000000000000011","111111111111111101","111111111111011100","000000000000101000","111111111111011001","000000000000010000","000000000000010100","111111111111111011","000000000000010010","111111111111101100","111111111111110111","000000000000011010","000000000000010100","111111111111111010","000000000000011111","000000000000100000","111111111111110000","000000000000101100","111111111111110110","111111111111110011","111111111111100100","000000000000101111","000000000000010100","000000000000000000","000000000000001001","111111111111110000","000000000000110000","000000000000100101","111111111111110111","111111111111111010","111111111111011110","111111111111111111","111111111111110000","000000000000001110","000000000000000010","000000000000000000","111111111111101001","111111111111101111","111111111111100111","111111111111110001","111111111111100001","111111111111110101","111111111111011110","111111111111110111","000000000000010100","111111111111101110","000000000000011100","111111111111111110","000000000000110101","111111111111101000","000000000000110100","000000000000101011","111111111111011001","000000000000001011","111111111111111110","111111111111110111","111111111111111100","000000000000000011","000000000000000001","000000000000010110","111111111111111110","000000000000000000","000000000000001010","000000000000100011","000000000000001011","111111111111011111","111111111111111010","111111111111110011","111111111111111101","000000000000000000","000000000000001011","111111111111110111","000000000000001010","000000000000000011","111111111111110010","000000000000010010","111111111111101111","000000000000001000","111111111111110001","000000000000101100","000000000000010000","000000000000001001","000000000000000000","000000000000100010","000000000000011111","000000000000000000","000000000000000000","000000000000001110","000000000000010110","111111111111110010","000000000000001011","111111111111110101","000000000000001010","000000000000011111","000000000000011110","000000000000000100","000000000000001111","111111111111011111","000000000000011000","000000000000000111","111111111111011111","111111111111111111","000000000000000000","111111111111100110","000000000000001010","111111111111011010","111111111111110100","111111111111110110"),
("000000000000001110","111111111111100011","000000000000000010","111111111111111010","111111111111110111","000000000000000010","000000000000100010","000000000000101010","000000000000100010","111111111111101010","111111111111101000","111111111111110000","000000000000001100","000000000000010100","000000000000000010","111111111111101000","000000000000000110","111111111111111100","000000000000001101","111111111111110000","111111111111100011","111111111111010110","111111111111101111","000000000000010101","111111111111101001","000000000000100001","000000000000011101","000000000000000100","000000000000101000","111111111111101001","111111111111111011","000000000000000011","111111111111110011","111111111111101100","000000000000011011","000000000000011110","111111111111111011","000000000000000011","111111111111111000","000000000000001001","111111111111111011","111111111111110100","111111111111110010","111111111111111000","000000000000000001","000000000000001100","000000000000000010","000000000000101100","111111111111110110","111111111111111011","111111111111110001","111111111111111010","111111111111100010","000000000000000011","000000000000101011","000000000000010011","000000000000000010","000000000000000111","111111111111101101","111111111111111110","111111111111110010","111111111111111110","000000000000000111","000000000000000010","000000000000001001","111111111111110111","000000000000001001","111111111111111001","000000000000011001","111111111111110110","000000000000000000","000000000000010010","111111111111100001","000000000000010110","111111111111110101","111111111111110100","111111111111110101","000000000000000110","000000000000000110","000000000000011100","000000000000000000","000000000000001001","000000000000001110","000000000000011001","000000000000000010","000000000000001001","000000000000000100","000000000000000101","000000000000100000","000000000000001110","000000000000001110","111111111111110111","111111111111111101","111111111111010111","000000000000000100","000000000000001011","111111111111101100","000000000000100010","111111111111100010","000000000000100000","000000000000011010","000000000000000001","111111111111110000","111111111111101000","111111111111111101","111111111111110001","000000000000001110","000000000000110000","000000000000011100","000000000000010001","111111111111110101","111111111111011100","000000000000100001","000000000000000111","000000000000101111","000000000000010100","000000000000001111","111111111111101010","000000000000001001","111111111111101100","111111111111101100","111111111111100000","000000000000011000","111111111111111001","000000000000011011","111111111111111110","111111111111110101","000000000000000100"),
("000000000000000001","111111111111100100","000000000000000110","000000000000000111","000000000000011111","000000000000100100","111111111111111111","000000000000101011","000000000000001111","111111111111100101","111111111111010101","111111111111100110","111111111111111011","111111111111111100","000000000000011010","111111111111110101","111111111111111011","111111111111110001","111111111111101111","111111111111111101","111111111111111100","111111111111011000","111111111111101101","000000000000000000","111111111111101110","111111111111111111","000000000000010001","000000000000010011","000000000000000101","000000000000000110","111111111111111000","000000000000010000","111111111111101111","111111111111111001","000000000000001011","000000000000000000","000000000000010001","000000000000001101","111111111111111010","111111111111110101","111111111111101101","111111111111011011","111111111111111101","000000000000011001","000000000000001000","000000000000100010","111111111111100010","000000000000101100","111111111111101101","111111111111101011","000000000000011001","000000000000000100","111111111111101011","111111111111110001","000000000000000000","000000000000010100","000000000000010101","000000000000000011","111111111111100000","000000000000010000","111111111111110010","000000000000001111","000000000000000010","000000000000010110","000000000000111000","111111111111111111","000000000000000001","000000000000000110","000000000000001101","111111111111100000","000000000000010111","111111111111101000","111111111111011101","000000000000101010","000000000000000011","000000000000000101","000000000000010011","111111111111111100","000000000000001010","000000000000000111","111111111111111000","111111111111111001","000000000000100101","000000000000010101","111111111111100011","000000000000011100","000000000000000001","000000000000010000","000000000000010111","111111111111110011","000000000000011001","111111111111110011","111111111111101101","111111111111111000","000000000000010000","000000000000001011","000000000000001011","000000000000000111","111111111111111100","111111111111111101","000000000000000100","111111111111101111","111111111111101100","111111111111111110","111111111111100100","000000000000001101","000000000000001101","000000000000010100","000000000000101110","000000000000001001","000000000000001001","111111111111001001","000000000000000100","000000000000010001","111111111111111100","000000000000010010","000000000000001010","000000000000000000","000000000000001010","111111111111111111","111111111111011111","111111111111111001","000000000000010111","000000000000001001","000000000000101011","111111111111101101","111111111111111011","000000000000100100"),
("000000000000000110","111111111111110001","000000000000100011","000000000000000101","111111111111111110","000000000000001101","000000000000010110","000000000000001011","111111111111111101","111111111111100001","111111111111001101","111111111111111000","000000000000000011","000000000000010100","000000000000101010","111111111111011100","000000000000001110","000000000000000011","111111111111111111","111111111111111111","111111111111111011","111111111111101111","111111111111111011","111111111111110011","000000000000000001","111111111111111111","000000000000010100","000000000000001110","111111111111110100","111111111111110111","000000000000000100","000000000000000110","000000000000000111","000000000000000101","111111111111111010","111111111111100000","000000000000011011","111111111111101110","000000000000000101","111111111111110101","111111111111011001","111111111111100111","111111111111111100","111111111111110010","000000000000011110","000000000000100101","111111111111101110","000000000000010011","000000000000010001","111111111111111000","000000000000010101","000000000000000110","111111111111111110","000000000000000010","000000000000001111","000000000000010101","000000000000011110","000000000000000100","000000000000100101","111111111111101010","000000000000001110","000000000000010101","111111111111111011","111111111111111000","111111111111110111","000000000000100110","111111111111011111","111111111111100110","111111111111111001","111111111111111100","111111111111110101","000000000000001000","000000000000000000","000000000000100011","111111111111111010","111111111111111101","000000000000001000","111111111111101110","000000000000010100","111111111111111100","000000000000001101","111111111111111111","000000000000011101","000000000000001101","111111111111101110","000000000001000001","000000000000001000","000000000000000000","111111111111111010","000000000000000010","000000000000010110","111111111111110111","111111111111100000","000000000000001001","000000000000101100","111111111111111100","000000000000000110","000000000000100010","000000000000010001","000000000000000011","111111111111110100","000000000000010001","111111111111101100","111111111111011010","111111111111110101","111111111111111001","000000000000010011","111111111111111111","000000000000101001","000000000000110101","000000000000010100","111111111111011100","000000000000001101","111111111111101101","000000000000001110","111111111111110000","111111111111110110","111111111111110111","111111111111101011","111111111111111101","111111111111110101","111111111111101011","000000000000010011","000000000000010000","000000000000010010","111111111111111111","000000000000000010","000000000000011001"),
("111111111111111100","111111111111110010","000000000000010000","111111111111101010","111111111111101110","000000000000000011","000000000000010011","111111111111111011","111111111111111100","111111111111101000","111111111111011110","111111111111110101","000000000000000100","000000000000001111","000000000000010000","111111111111011011","000000000000000110","111111111111101000","111111111111111000","111111111111101110","000000000000010010","111111111111110100","000000000000000000","111111111111110101","000000000000001111","111111111111110111","000000000000010110","111111111111111111","000000000000001000","000000000000001100","000000000000000011","000000000000000111","000000000000010110","000000000000010100","111111111111100001","111111111111100001","000000000000010101","111111111111100111","000000000000011000","000000000000010001","111111111111101100","000000000000001101","000000000000001000","111111111111101000","111111111111111001","000000000000000000","111111111111111010","000000000000000011","000000000000010111","111111111111110111","000000000000010101","000000000000001001","111111111111111001","111111111111111101","000000000000000100","000000000000001010","000000000000100001","000000000000001111","000000000000011011","111111111111101111","000000000000001011","111111111111110101","111111111111101100","000000000000001100","111111111111010111","000000000000010110","111111111111101010","111111111111111100","000000000000001111","000000000000000110","111111111111111110","111111111111110100","000000000000000101","000000000000000111","000000000000010010","000000000000000111","111111111111111100","111111111111111111","000000000000001011","000000000000011010","111111111111101110","111111111111111111","000000000000011010","000000000000011011","111111111111111010","000000000000101011","000000000000110000","111111111111100111","000000000000000001","000000000000000011","000000000000000101","000000000000001000","111111111111101101","111111111111101110","000000000000100100","000000000000000100","000000000000000000","000000000000111100","000000000000110001","111111111111101001","111111111111110000","000000000000000011","111111111111110000","111111111111011110","111111111111110000","111111111111110001","000000000000000001","000000000000011000","000000000000011101","000000000000010110","000000000000010011","000000000000001001","111111111111101011","000000000000001000","111111111111110100","000000000000011000","000000000000010001","000000000000000010","111111111111110111","111111111111110111","111111111111111010","000000000000000011","111111111111101000","111111111111101010","000000000000010000","000000000000000000","111111111111110110","000000000000001010"),
("111111111111101010","111111111111110010","111111111111110011","111111111111100010","000000000000000110","111111111111110111","000000000000011110","111111111111101011","111111111111111111","111111111111110001","111111111111000100","111111111111110101","111111111111101011","111111111111111010","000000000000100001","111111111111010000","000000000000001101","111111111111110001","111111111111111110","111111111111110010","000000000000000000","000000000000000101","111111111111111001","111111111111100011","111111111111101101","111111111111101110","000000000000001011","111111111111110101","000000000000100010","111111111111011010","111111111111101111","111111111111111110","111111111111111011","000000000000010111","111111111111111000","111111111111101111","111111111111101111","111111111111111011","111111111111111010","000000000000010101","000000000000001010","111111111111110100","111111111111111110","111111111111100100","000000000000011000","111111111111110000","000000000000011101","111111111111110101","111111111111111110","000000000000001010","000000000000011011","111111111111111010","111111111111111010","000000000000000011","111111111111011011","000000000000101000","000000000000000100","000000000000010111","000000000000000100","000000000000000111","000000000000000011","000000000000001000","000000000000000001","000000000000000111","111111111110011100","000000000000011001","111111111111101001","111111111111110001","000000000000010001","111111111111011010","000000000000001011","111111111111111100","000000000000000001","000000000000000010","000000000000001101","000000000000001110","000000000000000000","111111111111101101","000000000000101010","000000000000011111","111111111111101110","000000000000010010","000000000000001110","000000000000010011","111111111111100011","000000000000100111","000000000000001110","000000000000010111","000000000000000000","111111111111111011","000000000000000100","111111111111110110","111111111111110010","111111111111110101","000000000000000000","111111111111111010","000000000000000111","000000000000101100","000000000000100010","000000000000001110","000000000000010001","000000000000001001","111111111111101111","111111111111101000","000000000000000000","111111111111111101","111111111111111101","000000000000010101","111111111111101110","000000000000001001","111111111111110111","000000000000010100","111111111111110100","000000000000000111","111111111111110011","111111111111110111","111111111111111111","000000000000001011","111111111111011110","111111111111110101","111111111111110011","111111111111110110","111111111111111000","111111111111110100","000000000000011010","000000000000001111","111111111111101110","000000000000001001"),
("111111111111100001","000000000000001000","000000000000000000","111111111111110001","000000000000010001","111111111111100000","000000000000100111","000000000000011011","111111111111100101","111111111111110111","111111111111100101","111111111111110001","111111111111100111","111111111111110101","000000000000110000","111111111111101100","000000000000001000","111111111111110011","111111111111101011","111111111111011001","000000000000000100","000000000000101101","000000000000001010","111111111111101010","000000000000010001","000000000000000111","111111111111100001","111111111111101101","000000000000000011","111111111111101101","111111111111111100","000000000000010010","000000000000010000","000000000000001011","111111111111101100","111111111111110000","000000000000000110","000000000000000010","000000000000000000","000000000000011111","111111111111111111","111111111111110011","000000000000011000","111111111111100101","000000000000001000","000000000000000110","111111111111101100","111111111111111101","000000000000011111","000000000000010101","000000000000001001","000000000000000001","000000000000010100","000000000000000001","111111111111100101","000000000000001001","111111111111110101","000000000000010010","000000000000001100","111111111111111101","000000000000011000","111111111111111101","111111111111010001","111111111111111110","111111111111011001","111111111111111110","111111111111101101","111111111111110010","000000000000010110","111111111111101111","000000000000000111","111111111111101111","000000000000011111","111111111111111111","000000000000000000","000000000000011100","111111111111110000","111111111111110010","000000000000100100","000000000000000111","111111111111101010","000000000000000010","000000000000001110","000000000000010101","111111111111111100","000000000000001100","000000000000010001","000000000000010000","000000000000001110","000000000000011010","000000000000000011","000000000000010101","111111111111101010","000000000000011010","111111111111110111","111111111111110111","000000000000000010","000000000000011011","000000000000011000","000000000000001111","000000000000000011","111111111111101100","000000000000000000","111111111111100111","111111111111011110","111111111111101101","111111111111111000","000000000000010101","111111111111111000","000000000000000111","111111111111110011","000000000000100111","000000000000010100","000000000000011010","111111111111111100","000000000000010011","111111111111111111","111111111111101010","111111111111111110","000000000000011010","000000000000000110","111111111111111011","111111111111011100","000000000000000101","000000000000001111","000000000000000111","111111111111101110","111111111111110011"),
("111111111111110100","000000000000011000","000000000000010101","111111111111100111","111111111111110110","111111111111111100","000000000000100000","111111111111110001","000000000000000010","000000000000010101","111111111111100010","000000000000000011","111111111111101011","111111111111111010","000000000000010000","000000000000001011","000000000000010000","111111111111100100","111111111111110000","000000000000001101","000000000000000001","000000000000010100","111111111111111111","111111111111110111","111111111111111101","111111111111111001","000000000000000110","111111111111110001","000000000000010111","111111111111101010","111111111111011111","000000000000001110","111111111111110110","000000000000000010","000000000000001001","111111111111101110","111111111111111001","000000000000010010","000000000000000000","000000000000100000","000000000000010101","111111111111111111","000000000000001010","111111111111100001","111111111111101000","000000000000001110","111111111111101001","111111111111111001","000000000000000010","111111111111111001","000000000000011111","111111111111111101","000000000000001110","000000000000011001","111111111111110101","111111111111110000","111111111111101011","111111111111110110","111111111111111111","111111111111101101","000000000000000110","111111111111110000","111111111111111001","000000000000000010","000000000000001010","111111111111110100","111111111111010111","111111111111111000","000000000000100101","111111111111110001","111111111111100100","111111111111101101","111111111111101000","000000000000000010","000000000000100000","000000000000001111","111111111111110110","000000000000011000","000000000000001101","111111111111111010","111111111111111110","111111111111011110","000000000000011000","000000000000011100","111111111111100111","111111111111110011","000000000000001111","000000000000011010","000000000000000111","000000000000011000","111111111111101111","111111111111111010","111111111111111100","000000000000000111","000000000000000000","111111111111011101","000000000000001111","000000000000100111","000000000000010100","111111111111110100","000000000000000011","000000000000000101","111111111111111111","111111111111001110","000000000000000011","000000000000001000","111111111111100011","000000000000001000","111111111111011100","000000000000010001","111111111111101100","000000000000001010","111111111111111001","000000000000010111","111111111111111001","000000000000010100","000000000000000001","111111111111110101","111111111111100010","000000000000010101","000000000000010100","111111111111111101","111111111111111011","111111111111010001","000000000000001110","000000000000010110","111111111111110110","111111111111101010"),
("111111111111001101","000000000000011110","000000000000001100","111111111111111001","000000000000010000","000000000000000010","000000000000000011","000000000000000101","000000000000010011","000000000000000100","111111111111011001","000000000000000010","111111111111010010","111111111111101001","000000000000100100","111111111111101110","000000000000000000","111111111111100110","111111111111101111","000000000000001000","111111111111110011","000000000000001101","111111111111111111","000000000000000000","111111111111101000","000000000000000011","111111111111101011","111111111111101011","000000000000001100","111111111111100000","111111111111101111","000000000000010100","000000000000001100","111111111111110011","000000000000001010","111111111111110100","111111111111111010","000000000000000011","111111111111011011","000000000000100000","000000000000001101","000000000000010000","000000000000000010","111111111111010011","111111111111110001","000000000000101110","000000000000011001","000000000000001101","000000000000001101","000000000000001001","000000000000011001","111111111111100100","111111111111111010","000000000000001101","000000000000000101","000000000000001110","111111111111111010","000000000000010110","000000000000001111","000000000000001010","111111111111111110","111111111111101110","111111111111101010","000000000000010101","000000000000000110","111111111111111111","111111111111001001","000000000000010100","000000000000110110","000000000000000101","111111111111101011","111111111111011000","111111111111100000","000000000000010111","000000000000000101","000000000000110010","111111111111100110","111111111111110101","000000000000010110","000000000000100011","000000000000000111","111111111111011011","000000000000010110","111111111111100010","111111111111100000","000000000000001000","000000000000011101","000000000000100001","111111111111111111","000000000000101100","000000000000000100","000000000000000010","000000000000010011","000000000000000010","111111111111111001","111111111111101001","000000000000010010","000000000000011011","111111111111110111","000000000000000110","111111111111110110","111111111111110100","000000000000011010","111111111111100001","111111111111011111","000000000000000101","000000000000000001","000000000000011011","111111111111001101","000000000000000101","111111111111111000","000000000000000100","000000000000001000","000000000000010101","111111111111101011","000000000000001100","000000000000010010","000000000000000010","111111111111011111","000000000000100011","111111111111101011","111111111111110100","111111111111100111","111111111111100100","000000000000001100","111111111111111101","111111111111101100","111111111111111101"),
("111111111111110111","000000000000010011","000000000000010110","111111111111001100","000000000000000100","111111111111110011","111111111111111100","000000000000010001","111111111111111100","000000000000001000","111111111111110001","000000000000110011","111111111111010111","111111111111001110","000000000000001010","111111111111110110","000000000000010011","111111111111101011","000000000000000011","000000000000001001","000000000000001001","000000000000100011","000000000000010000","111111111111101000","000000000000001111","111111111111110010","000000000000000111","111111111111111011","000000000000001001","111111111111110011","111111111111110011","111111111111111101","000000000000001101","111111111111100111","000000000000001010","111111111111100001","111111111111111111","111111111111110000","111111111111001111","000000000000010100","000000000000101100","111111111111110001","000000000000001011","111111111111101111","111111111111101100","000000000000010010","000000000000011010","111111111111111110","000000000000010111","111111111111110111","000000000000010001","000000000000001010","000000000000010111","111111111111111010","000000000000010100","111111111111111011","111111111111011100","000000000000000010","000000000000000000","000000000000010010","000000000000010001","111111111111101100","111111111111110110","111111111111110101","111111111111110101","000000000000001101","111111111111011010","000000000000000101","000000000000111010","000000000000011001","111111111111101110","111111111111011010","111111111111100010","000000000000001010","000000000000000110","000000000000011111","111111111111101101","111111111111101010","111111111111111100","000000000000000000","000000000000000000","111111111111001101","000000000000000000","111111111111001110","000000000000000010","000000000000000111","000000000000110000","000000000000011101","000000000000000000","000000000000001110","000000000000010000","000000000000000000","000000000000100100","000000000000001000","111111111111110101","111111111111011111","000000000000100101","111111111111110101","111111111111011000","000000000000000100","111111111111100101","000000000000001000","111111111111111111","111111111111011001","111111111111111001","000000000000011000","111111111111101010","000000000000001101","111111111111100010","111111111111101000","111111111111100100","111111111111110010","000000000000001100","000000000000010110","111111111111101001","000000000000001110","000000000000010001","111111111111101101","111111111111100101","000000000000011000","111111111111011100","111111111111111011","111111111111111001","111111111111001101","000000000000101100","000000000000010110","000000000000001101","000000000000010001"),
("111111111111111011","000000000000010010","111111111111111010","111111111111110100","111111111111111111","111111111111110001","000000000000000100","000000000000010111","111111111111111001","000000000000101100","000000000000001010","000000000000100010","000000000000000000","111111111111100000","111111111111010000","000000000000101110","111111111111111010","111111111111110011","111111111111110010","000000000000011001","000000000000101111","111111111111110001","000000000000001001","111111111111110011","000000000000001000","111111111111110100","111111111111101011","111111111111101100","111111111111110101","000000000000010110","000000000000001011","111111111111110110","000000000000010100","111111111111100110","111111111111101110","000000000000001100","000000000000001010","111111111111111000","111111111111100111","111111111111111111","000000000000011101","111111111111111110","000000000000100110","111111111111111111","000000000000000000","111111111111100001","000000000000101100","000000000000001111","111111111111101110","111111111111011000","000000000000110100","000000000000010001","000000000000000000","111111111111100000","000000000000000010","111111111111100110","111111111111100010","000000000000010001","111111111111100100","000000000000010000","111111111111111110","000000000000000000","111111111111110111","111111111111101101","111111111111111001","111111111111111101","111111111111001011","000000000000010010","000000000000110100","111111111111111110","000000000000001010","111111111111101011","111111111111011011","000000000000001100","111111111111110111","000000000000100110","111111111111101001","111111111111100011","111111111111001001","000000000000011110","111111111111110101","111111111111010010","000000000000001101","111111111111100111","000000000000000111","111111111111011011","000000000000011110","000000000000100010","111111111111000110","111111111111110001","111111111111111011","000000000000000000","000000000000000100","000000000000011000","000000000000000011","111111111111111011","000000000000110001","000000000000001010","111111111111100111","111111111111100100","000000000000001000","111111111111110000","111111111111101011","111111111111101000","111111111111111110","000000000000100011","111111111111110001","111111111111110111","111111111111011110","111111111111110100","111111111111100010","111111111111111111","000000000000000101","111111111111110100","000000000000000000","000000000000000001","000000000000000101","000000000000100000","111111111111101000","000000000000011000","111111111111101101","000000000000001111","111111111111110000","111111111111011001","000000000000010111","111111111111111111","000000000000101101","111111111111100101"),
("000000000000100000","000000000000100011","111111111111110110","111111111111111001","000000000000000010","000000000000100110","000000000000010111","000000000000010011","000000000000001101","111111111111110011","111111111111111111","000000000000010010","111111111111100001","111111111110110100","111111111111110101","000000000000011001","111111111111110010","000000000000001101","111111111111011001","111111111111111000","000000000000000000","111111111111110000","000000000000001100","000000000000000011","000000000000000000","000000000000001100","111111111111010001","111111111111101000","111111111111110010","111111111111101111","111111111111111011","000000000000000111","000000000000010010","111111111111101110","000000000000000000","000000000000001000","000000000000001000","111111111111110100","111111111111001110","111111111111101001","111111111111101111","111111111111101001","000000000000111001","000000000000101011","000000000000000101","111111111111011110","000000000000001001","000000000000110000","111111111111011111","111111111111101010","000000000000000010","111111111111111010","111111111111111101","111111111111001011","000000000000001100","111111111111111101","111111111111111010","111111111111110100","111111111111101111","000000000000001001","111111111111001101","111111111111111111","111111111111101110","000000000000001011","111111111111110011","111111111111101010","111111111111110001","000000000000101101","111111111111101111","111111111111011101","000000000000001111","111111111111011011","111111111110111101","000000000000001111","000000000000000001","000000000000001110","000000000000100110","111111111111110100","111111111111101010","000000000000010100","111111111111101100","000000000000001100","000000000000111100","111111111111010000","111111111111110110","111111111111011010","111111111111011111","000000000000001101","000000000000000001","111111111110110101","111111111111110111","111111111111101110","000000000000001101","000000000000010100","111111111111110011","111111111111111100","000000000000100111","000000000000000101","111111111111100010","111111111111111011","000000000001000001","111111111111110100","111111111111010111","111111111111110101","111111111111101010","000000000000100101","111111111111101000","111111111111110111","111111111111101111","000000000000000110","111111111111100110","111111111111100111","000000000000011001","111111111111111000","111111111110110111","000000000000000001","000000000000011101","000000000000000000","111111111111010110","111111111111110101","000000000000000011","000000000001010011","000000000000001110","000000000000011011","000000000000011111","000000000000000110","000000000000011110","000000000000000011"),
("111111111111111010","111111111111101000","111111111111110100","000000000000001000","000000000000010100","000000000000110110","000000000000010010","000000000000001011","000000000000010111","111111111111000000","000000000000010100","111111111111100111","000000000000001100","111111111111111101","111111111111110001","111111111111110110","000000000000010001","111111111111101000","111111111111001110","000000000000101110","000000000000000110","111111111111101110","000000000000001011","111111111111011000","111111111111100100","000000000000001001","111111111111100100","111111111111111111","000000000000010001","000000000000000010","000000000000100110","111111111111100110","111111111111111110","111111111111010000","000000000000001000","111111111111110110","000000000000000000","000000000000101100","111111111111101100","000000000000011101","111111111111100001","111111111111110011","111111111111110111","111111111111111001","000000000000000000","111111111111111000","111111111111100000","000000000000011000","111111111111100111","111111111111111010","111111111111111111","000000000000011110","111111111111000001","111111111111111110","000000000000101100","000000000000101110","111111111111101010","000000000000001011","111111111111011101","000000000000001111","111111111111101100","000000000000010011","111111111111111110","000000000000000111","111111111111101010","111111111111001101","111111111111100011","111111111111011000","000000000000010110","111111111111101011","000000000000010011","000000000000010110","111111111111011101","000000000000010110","111111111111011100","000000000000001011","000000000000101111","000000000000001110","000000000000001001","000000000000101110","111111111111110001","000000000000011101","000000000001000111","000000000000000011","000000000000010010","111111111111101001","000000000000011111","000000000000101010","111111111111100001","111111111111100011","111111111111100100","111111111111011111","111111111111100010","111111111111111110","000000000000000000","000000000000011000","000000000000010101","000000000000011100","111111111111011100","000000000000011000","000000000000100101","111111111111110010","111111111111101001","000000000000000011","111111111111110100","000000000000011100","000000000000000000","111111111111011011","000000000000000001","111111111111110110","111111111111110010","000000000000011110","111111111111110111","111111111111110110","000000000000001000","111111111111111000","111111111111010101","000000000000010100","111111111111111011","000000000000011101","000000000000000101","000000000000100001","000000000000000100","000000000000001001","000000000000011001","111111111111011001","111111111111110011","000000000000000011"),
("000000000000101011","111111111111101101","111111111111011110","000000000000001110","111111111111101110","000000000000101001","000000000000001001","111111111111111111","111111111111111110","111111111111100011","000000000000001000","111111111111110111","000000000000001101","111111111111101100","111111111111100111","000000000000010011","000000000000101100","000000000000010101","111111111111110011","000000000000100111","000000000000100110","111111111111111100","000000000000000101","111111111111111101","111111111111011101","000000000000010111","000000000000001110","000000000000010001","000000000000010010","000000000000000110","000000000000010000","000000000000000111","000000000000000110","111111111111100000","000000000000001100","111111111111110011","000000000000001001","000000000000000100","111111111111110011","111111111111110010","000000000000000000","111111111111101011","000000000000101101","000000000000101010","111111111111111011","111111111111100001","111111111111110011","000000000000101110","111111111111101100","111111111111100101","111111111111111111","000000000000100000","111111111111011001","000000000000011010","000000000000001000","000000000000101000","111111111111101001","000000000000010010","111111111111001110","000000000000010001","111111111111110100","000000000000011011","000000000000100000","000000000000001110","111111111111111101","111111111111100100","111111111111111111","111111111111101110","000000000000001111","111111111111111001","000000000000011110","000000000000001100","111111111111111010","000000000000011000","000000000000000000","000000000000011001","000000000000001010","000000000000010000","111111111111110111","000000000000000011","000000000000000101","000000000000000000","000000000000100101","111111111111111001","000000000000000100","111111111111011110","111111111111110011","000000000000010110","111111111111111101","111111111111110110","111111111111110110","111111111111111100","111111111111110010","000000000000011011","111111111111011101","111111111111101010","000000000000010111","000000000000100011","111111111111100000","111111111111110101","000000000000001111","111111111111100100","111111111111101011","000000000000001100","111111111111110100","000000000000101100","111111111111100000","000000000000000001","000000000000001010","111111111111101101","111111111111110101","000000000000100010","000000000000001001","111111111111111101","000000000000010001","111111111111111100","111111111111101100","000000000000010100","111111111111111011","000000000000000000","000000000000001001","000000000000011001","000000000000001010","000000000000010101","000000000000101111","111111111111110101","000000000000011110","111111111111111000"),
("000000000000000111","000000000000001111","000000000000000001","000000000000000110","111111111111110001","000000000000000101","111111111111110001","111111111111101101","000000000000010000","000000000000001110","000000000000000000","111111111111110010","000000000000001100","111111111111110011","000000000000001100","111111111111111011","000000000000000101","111111111111111111","000000000000001001","111111111111110010","000000000000000000","000000000000000101","111111111111110100","111111111111101100","000000000000010000","000000000000001110","000000000000000010","111111111111110000","000000000000010101","000000000000001011","111111111111111111","000000000000001001","000000000000010001","111111111111110011","111111111111101111","000000000000001110","000000000000001101","000000000000001101","000000000000000010","111111111111111001","000000000000000000","111111111111110101","111111111111110010","111111111111110011","111111111111111101","111111111111101111","000000000000000011","000000000000000000","000000000000001110","111111111111111001","111111111111111000","000000000000000111","000000000000001000","111111111111101101","000000000000001001","000000000000001101","111111111111101110","000000000000000011","000000000000000110","000000000000001011","000000000000010010","000000000000000111","111111111111111110","111111111111110110","111111111111110011","111111111111111001","000000000000001001","111111111111111001","000000000000000000","000000000000001011","000000000000001000","000000000000000000","000000000000001011","000000000000001011","111111111111101010","000000000000010001","000000000000001000","111111111111110101","111111111111110001","000000000000000111","000000000000001011","000000000000010001","000000000000001110","111111111111110011","000000000000010001","111111111111110001","111111111111110100","111111111111111011","111111111111111111","111111111111111001","000000000000001011","111111111111110001","111111111111110111","111111111111101100","000000000000000100","000000000000010000","111111111111110111","111111111111111010","000000000000010001","111111111111110011","111111111111101110","111111111111111111","111111111111110100","111111111111101110","000000000000000000","111111111111110101","111111111111110011","000000000000001010","000000000000010011","000000000000000111","111111111111111000","111111111111110101","000000000000010001","111111111111110001","111111111111110110","111111111111101110","000000000000000010","000000000000001110","000000000000000111","111111111111110100","000000000000001010","000000000000000001","000000000000000000","000000000000001110","000000000000000000","111111111111110101","000000000000000001","000000000000001101"),
("000000000000000000","000000000000000010","000000000000001011","000000000000001110","000000000000000110","000000000000010000","111111111111110001","111111111111111000","000000000000000100","111111111111110111","000000000000000100","111111111111111011","111111111111110100","111111111111111111","000000000000001100","111111111111100000","000000000000000101","111111111111110111","000000000000001001","000000000000001001","111111111111101000","111111111111101100","000000000000001101","111111111111011110","111111111111101101","000000000000010010","000000000000000101","000000000000010100","000000000000011011","000000000000011100","111111111111011101","000000000000000100","000000000000010011","111111111111110110","111111111111100010","000000000000000110","111111111111110010","000000000000011010","000000000000000100","000000000000011111","000000000000010001","111111111111100011","000000000000010101","000000000000010010","000000000000001111","000000000000011011","111111111111111110","111111111111100111","000000000000010000","000000000000001001","000000000000011001","111111111111110111","000000000000000110","000000000000001110","000000000000001111","111111111111111100","111111111111111010","000000000000011111","111111111111110000","000000000000001110","111111111111111010","000000000000010010","000000000000000001","000000000000011101","000000000000000011","111111111111011001","111111111111011111","111111111111110100","000000000000000000","111111111111111001","000000000000001010","000000000000011110","111111111111110000","000000000000010110","000000000000100001","111111111111110011","000000000000000000","000000000000011110","111111111111111011","000000000000011000","000000000000010111","000000000000001010","111111111111101011","000000000000100000","000000000000010110","111111111111100110","111111111111100011","000000000000011111","000000000000001110","000000000000001101","000000000000000110","111111111111111001","000000000000010001","000000000000000101","111111111111111101","000000000000010101","000000000000000111","000000000000000101","000000000000010011","000000000000000010","111111111111100011","111111111111110101","000000000000000110","111111111111111101","111111111111111101","000000000000000110","000000000000010110","000000000000010001","000000000000000000","111111111111100111","111111111111111010","111111111111101010","000000000000010010","000000000000100001","000000000000000010","000000000000010101","000000000000011011","111111111111111101","000000000000000111","000000000000001011","000000000000000001","111111111111111100","111111111111101011","111111111111110111","111111111111101111","111111111111101011","111111111111111011","000000000000100011"),
("000000000000001110","000000000000011101","111111111111101010","111111111111110011","000000000000000011","000000000000000101","111111111111011111","000000000000101011","000000000000011010","111111111111110110","000000000000001100","000000000000101001","111111111111111001","000000000000000101","111111111111100110","111111111111110001","000000000000100000","111111111111111110","000000000000000011","000000000000001001","111111111111101010","111111111111110010","000000000000100100","000000000000000011","111111111111110101","111111111111111101","000000000000000111","111111111111110110","000000000000100001","000000000000010011","000000000000001010","000000000000000111","000000000000010001","000000000000001101","111111111111111101","000000000000000111","111111111111100001","000000000000100001","000000000000010110","000000000000000000","000000000000011111","111111111111111100","111111111111111111","000000000000010001","000000000000011001","111111111111110110","111111111111111101","111111111111110110","000000000000000100","111111111111110110","000000000000001111","000000000000011100","111111111111110100","000000000000000000","000000000000001010","111111111111100100","111111111111111101","000000000000000000","111111111111101010","000000000000000110","000000000000010011","000000000000001110","111111111111111110","000000000000010100","000000000000011111","111111111111010000","111111111111101100","000000000000000111","000000000000001100","111111111111111000","000000000000011001","000000000000010111","111111111111110110","000000000000001011","000000000000100100","000000000000000001","111111111111111000","111111111111110111","111111111111100100","000000000000011000","000000000000010001","111111111111101110","000000000000010000","111111111111110011","000000000000010001","000000000000001100","111111111111111001","000000000000100011","000000000000000001","111111111111110111","111111111111110111","111111111111111010","111111111111001001","111111111111110001","111111111111110101","111111111111110101","111111111111111011","111111111111101010","111111111111111011","000000000000010111","000000000000000101","111111111111110110","000000000000001011","000000000000011000","000000000000001110","000000000000000010","000000000000001011","111111111111100111","111111111111110001","111111111111110001","000000000000000010","111111111111110101","000000000000010000","000000000000010000","000000000000011001","000000000000001010","000000000000010100","000000000000000101","000000000000011010","000000000000011100","111111111111110101","111111111111101101","111111111111110100","000000000000110110","000000000000010111","111111111111101010","000000000000000011","111111111111111111"),
("000000000000001011","111111111111111110","111111111111100011","000000000000010110","000000000000010001","000000000000001111","111111111111100110","111111111111100101","000000000000000001","000000000000000000","111111111111001000","111111111111111111","111111111111101110","000000000000000000","111111111111110000","111111111111111111","000000000000110001","000000000000011011","000000000000011111","000000000000001111","111111111111110100","111111111111111101","111111111111110000","111111111111111100","111111111111111000","000000000000001101","111111111111111100","000000000000000000","000000000000011100","000000000000010001","000000000000110101","000000000000000000","000000000000011001","111111111111110111","000000000000010101","111111111111111101","000000000000010000","000000000000011011","111111111111100111","000000000000000001","111111111111110011","111111111111110111","000000000000011001","000000000000000101","000000000000010010","111111111111100110","111111111111111100","000000000000101001","111111111111101111","111111111111111010","000000000000010111","000000000000001100","111111111111110100","111111111111101101","000000000000101010","000000000000011011","111111111111011000","111111111111110000","111111111111000110","111111111111111110","111111111111100111","000000000000110000","000000000000010100","000000000000000100","111111111111110100","111111111111011101","111111111111101001","000000000000000011","111111111111100111","111111111111111100","111111111111111111","000000000000011001","111111111111100011","000000000000001001","111111111111111111","111111111111111000","111111111111111101","000000000000000010","111111111111101100","000000000000011010","111111111111011100","111111111111110110","000000000000000110","111111111111001010","000000000000000011","111111111111101001","000000000000100001","000000000000010100","000000000000000000","000000000000011010","000000000000000101","111111111111111000","111111111111110010","111111111111111000","000000000000000000","111111111111100101","000000000000010101","000000000000100110","111111111111110101","111111111111100110","000000000000001001","111111111111101111","111111111111101100","000000000000000111","111111111111101010","111111111111111110","111111111111011001","111111111111010110","111111111111100111","111111111111011010","111111111111111100","111111111111111101","000000000000001110","111111111111110101","000000000000011001","111111111111101111","111111111111111001","000000000000011011","111111111111011101","000000000000010110","111111111111110000","111111111111101100","111111111111111101","000000000000010011","000000000000011100","111111111111001001","111111111111100111","111111111111100010"),
("111111111111111110","111111111111111100","111111111111111111","111111111111111011","000000000000001100","000000000000000011","111111111111101011","000000000000001101","111111111111011101","000000000000000101","111111111110100011","111111111111010001","111111111111001011","111111111111100010","000000000000011001","000000000000000000","000000000000000011","000000000000000110","111111111111101111","000000000000100100","000000000000010000","000000000000000001","000000000000000111","111111111111111011","000000000000010001","111111111111111110","111111111111111011","000000000000000101","000000000000000101","000000000000010100","111111111111111111","000000000000000001","000000000000111010","111111111111110110","000000000000000001","111111111111000010","000000000000000000","111111111111101111","111111111111011100","000000000000010000","000000000000000001","111111111111010111","000000000000011001","111111111111101000","111111111111111110","111111111111110110","111111111111100011","000000000000001010","111111111111110011","000000000000001100","000000000000001110","000000000000000110","000000000000001011","111111111111110011","000000000000000100","000000000000010011","111111111111100010","000000000000010100","000000000000011000","111111111111111101","000000000000001111","000000000000110100","111111111111110101","111111111111110011","000000000000000100","000000000000000110","000000000000101010","111111111111110001","111111111111011100","000000000000001111","000000000000000101","000000000000000010","000000000000101110","000000000000000000","111111111111101100","111111111110110110","111111111111111010","000000000000011111","111111111111111011","111111111111111110","111111111111110101","000000000000010000","000000000000010101","000000000000001010","000000000000000110","111111111111101011","111111111111110110","000000000000001001","111111111111110101","000000000000010010","111111111111100011","111111111111111000","111111111111101101","000000000000000111","000000000000010110","000000000000001001","000000000000010010","000000000000000101","000000000000110000","000000000000001011","111111111111101111","111111111111011101","000000000000011100","111111111111100000","111111111111101101","000000000000010100","111111111111110011","111111111111101101","111111111111011101","111111111111101000","111111111111011111","000000000000001011","111111111111111010","000000000000010111","000000000000010101","000000000000000110","000000000000010111","111111111111101101","111111111111110111","000000000000000101","111111111111010011","111111111111100111","000000000000011101","111111111111101010","111111111111111000","111111111111011101","111111111111110110","000000000000001101"),
("000000000000010001","000000000000100010","000000000000100100","000000000000000111","000000000000001100","000000000000011010","111111111111110100","111111111111111100","111111111111100100","000000000000100000","111111111110011101","111111111111100001","111111111111100101","000000000000000111","000000000000010101","000000000000000011","000000000000100011","000000000000000011","111111111111100101","111111111111111011","000000000000011011","000000000000001100","000000000000011010","000000000000001010","000000000000000001","000000000000010010","111111111111011100","000000000000010001","000000000000000100","111111111111100010","000000000000011100","000000000000001001","000000000000010110","111111111111011011","111111111111111110","111111111111010100","111111111111110111","111111111111110100","111111111111111000","000000000000001111","111111111111110000","111111111111011001","111111111111111011","111111111111001100","000000000000001110","111111111111100010","111111111111111101","000000000000010101","111111111111111110","111111111111011101","000000000000011010","000000000000011101","000000000000000100","111111111111001010","111111111111100100","000000000000001010","111111111111011100","000000000000011000","111111111111110010","000000000000000010","000000000000001111","000000000001001011","111111111111111100","111111111111101110","111111111111101011","000000000000000110","000000000000010110","111111111111111010","111111111111011111","111111111111110011","111111111111110010","111111111111111110","000000000000111100","111111111111011010","111111111111110001","111111111111110001","111111111111111000","000000000000000100","000000000000000001","000000000000001100","111111111111111010","111111111111110110","000000000000000100","111111111111100111","000000000000000001","111111111111101011","111111111111100000","000000000000001111","111111111111101010","000000000000000001","111111111111111001","000000000000000111","000000000000000010","000000000000100010","111111111111110110","111111111111101010","000000000000000110","000000000000001101","000000000000010111","000000000000000001","000000000000011011","111111111111110101","000000000000001011","111111111111100011","111111111111101101","000000000000010000","111111111111011110","111111111111111001","111111111111100000","000000000000001110","111111111111110000","000000000000000000","000000000000000101","000000000000000101","111111111111110001","000000000000010010","000000000000000111","111111111111011100","111111111111101110","111111111111101101","111111111111011110","111111111111011110","111111111111110010","111111111111110011","111111111111110100","111111111111111001","000000000000000100","111111111111011001"),
("000000000000100110","000000000000110101","000000000000100010","111111111111110110","111111111111111011","000000000000010101","000000000000000100","111111111111101010","111111111111011011","111111111111111000","111111111110100000","111111111111101010","000000000000010010","000000000000001001","000000000000101000","000000000000001001","000000000000000000","000000000000000000","111111111111011111","000000000000000011","111111111111110111","000000000000100110","000000000000000010","000000000000010000","000000000000010010","000000000000000001","111111111111101110","111111111111101001","000000000000000001","111111111111010111","000000000000000100","111111111111111011","111111111111111000","111111111111101010","111111111111011111","111111111111100000","000000000000010000","000000000000000111","111111111111101010","000000000000000000","111111111111010100","111111111111101011","111111111111110111","111111111111000111","111111111111110111","111111111111100011","000000000000001010","000000000000011110","111111111111100111","111111111111111101","000000000000000000","000000000000100000","000000000000001010","111111111111100111","111111111111100010","000000000000010010","111111111111010001","000000000000000000","000000000000000010","000000000000000110","111111111111110110","000000000000101100","000000000000011000","111111111111110110","111111111111100000","000000000000001110","000000000000100011","111111111111111111","000000000000011010","000000000000000011","111111111111110111","111111111111110111","000000000000010001","111111111111111111","111111111111101110","111111111111000111","000000000000100010","111111111111110000","000000000000010111","000000000000010111","111111111111101100","111111111111101111","000000000000100111","111111111111101010","111111111111110001","111111111111110111","111111111111011101","111111111111110100","111111111111110000","000000000000000010","000000000000001010","111111111111110010","111111111111111000","000000000000000101","000000000000000101","111111111111001110","111111111111011111","000000000000001010","111111111111101101","000000000000001000","000000000000000100","000000000000000101","111111111111110000","000000000000000101","111111111111111010","000000000000010101","111111111111111101","000000000000010101","111111111111010110","000000000000000110","000000000000001001","111111111111110000","000000000000010100","111111111111110110","000000000000010011","000000000000010001","000000000000001110","111111111111010000","111111111111010011","111111111111010100","111111111111110100","111111111111100100","111111111111101101","000000000000000111","000000000000011000","111111111111111100","111111111111110001","111111111111111000"),
("000000000000010011","000000000000111011","000000000000001100","111111111111110101","000000000000011001","000000000000011000","000000000000010110","000000000000000011","111111111111101110","000000000000100011","111111111110010100","111111111111111000","111111111111111000","000000000000000000","000000000000001101","111111111111111100","000000000000100001","111111111111111111","111111111110111010","000000000000010110","000000000000001001","000000000000110010","000000000000011011","000000000000001000","111111111111111110","000000000000000111","111111111111101110","000000000000000000","000000000000001001","111111111111100001","000000000000001001","111111111111110111","111111111111111001","111111111111110010","111111111111100110","111111111111110010","000000000000000110","111111111111101101","111111111111100011","000000000000000000","111111111111101011","111111111111011011","111111111111110001","111111111111010001","111111111111111000","000000000000001011","111111111111101000","000000000000011011","111111111111101101","000000000000001101","000000000000001101","000000000000000011","000000000000011101","111111111111010011","111111111110111100","000000000000000001","111111111111100111","000000000000001101","000000000000011001","111111111111111011","111111111111111000","000000000000010001","000000000000010110","000000000000100011","111111111111001000","000000000000010001","000000000000000000","000000000000000000","000000000000110011","000000000000010011","111111111111111010","111111111111111001","000000000000011111","000000000000011100","111111111111111110","111111111111011111","000000000000000111","111111111111110100","000000000000100011","000000000000101101","000000000000001010","111111111111101110","000000000000100111","000000000000000000","111111111111011111","000000000000000000","111111111111011100","111111111111111101","000000000000000000","111111111111101111","000000000000011010","111111111111111000","111111111111101100","000000000000000100","111111111111110011","111111111111100100","111111111111101101","111111111111110110","111111111111100011","111111111111100111","000000000000011000","111111111111101111","111111111111110111","111111111111101011","111111111111110111","000000000000011001","111111111111110110","000000000000000001","111111111111100101","000000000000011101","111111111111111111","111111111111100011","000000000000000011","111111111111101000","000000000000001101","111111111111111010","111111111111110111","111111111111000011","111111111111010111","111111111111010111","111111111111110010","111111111111100001","111111111111100101","111111111111110101","000000000000100001","111111111111101010","111111111111111001","111111111111111101"),
("000000000000010011","000000000000101001","000000000000110001","111111111111111100","111111111111111111","000000000000100101","000000000000011110","111111111111111111","111111111111111001","111111111111111110","111111111110001101","000000000000010000","111111111111100100","000000000001000111","000000000000001000","000000000000010000","000000000000001110","111111111111111000","111111111111001010","111111111111111111","000000000000010000","000000000000010000","000000000000000101","000000000000011000","000000000000001011","111111111111101111","000000000000000000","111111111111011101","000000000000100010","000000000000000101","000000000000001011","111111111111110111","111111111111100110","111111111111111110","111111111111010101","111111111111010001","000000000000000011","111111111111101111","111111111111110110","111111111111100011","111111111111100000","111111111111111111","111111111111101001","000000000000001101","111111111111111111","000000000000010110","111111111111010100","000000000000110111","000000000000001110","000000000000001111","000000000000110010","000000000000000011","000000000000000010","111111111111100100","111111111111010000","000000000000100010","111111111111101011","111111111111101010","000000000000100101","111111111111111010","000000000000001000","000000000000000010","000000000000010011","000000000000001110","111111111111010110","000000000000101011","111111111111111111","111111111111100101","000000000001001001","000000000000010111","000000000000001001","111111111111101101","000000000000000011","111111111111110101","111111111111100100","111111111110111000","000000000000011001","111111111111110111","000000000000010010","000000000000011101","000000000000011101","111111111111100000","000000000000001000","111111111111111101","111111111111101111","000000000000011000","111111111111011110","111111111111101101","000000000000011011","000000000000011000","000000000000001100","111111111111101101","000000000000000110","000000000000010010","111111111111100101","111111111111111010","111111111111101100","111111111111111001","111111111111011100","111111111111111111","000000000000000101","111111111111111000","000000000000000110","111111111111100010","111111111111100111","000000000000000010","000000000000001100","111111111111101001","111111111111100000","000000000000010010","000000000000001010","000000000000000000","000000000000000000","111111111111100001","111111111111111011","000000000000011001","000000000000001001","111111111111010001","111111111111010110","111111111111000111","000000000000000010","111111111111110011","111111111111101100","111111111111000000","000000000000010101","111111111111100111","111111111111111101","111111111111110000"),
("000000000000010111","000000000000010110","000000000000101100","000000000000000011","000000000000011000","000000000000000000","000000000000011101","000000000000001101","111111111111111101","000000000000010001","111111111111000100","000000000000000001","111111111111100111","000000000000101000","111111111111101100","000000000000011010","000000000000010001","111111111111110111","111111111111011111","000000000000000001","111111111111110011","111111111111100100","000000000000001001","111111111111110010","000000000000000010","000000000000000001","111111111111100010","111111111111111010","000000000000010011","111111111111111001","000000000000000000","000000000000000010","111111111111101101","111111111111010111","111111111111100001","111111111111100110","000000000000000100","111111111111100101","000000000000001100","111111111111101111","111111111111010010","111111111111111100","111111111111110010","000000000000000101","000000000000010010","000000000000001011","111111111111101001","000000000000010110","111111111111101011","000000000000000100","000000000000101010","000000000000001011","000000000000100001","111111111111011000","111111111110111000","000000000000000000","111111111111011001","111111111111111100","000000000000001001","111111111111111101","111111111111101010","111111111111111000","000000000000001111","000000000000011000","111111111111001110","000000000000010001","111111111111101110","000000000000001010","000000000001001011","111111111111110100","000000000000010100","111111111111101100","111111111111110101","111111111111101110","111111111111110111","111111111111001101","000000000000011001","000000000000001000","000000000000010111","000000000000001001","000000000000000011","111111111111110110","000000000000011001","000000000000001111","000000000000000011","000000000000001001","111111111111110100","111111111111110111","000000000000100001","000000000000100001","000000000000010111","111111111111110111","000000000000000101","000000000000001111","111111111111100111","111111111111100101","111111111111110010","000000000000000010","111111111111000110","111111111111110110","000000000000101001","111111111111111111","000000000000001100","000000000000000000","000000000000001111","000000000000101001","000000000000010101","111111111111010101","111111111111111010","000000000000001001","000000000000010101","111111111111110100","000000000000011101","111111111111110100","000000000000010100","000000000000010111","000000000000000011","111111111111010100","111111111111010111","111111111111101000","000000000000001010","000000000000001111","111111111111010001","111111111110111010","000000000000011000","111111111111101111","000000000000010101","111111111111110101"),
("000000000000010110","111111111111111010","000000000000101001","000000000000000000","111111111111101101","000000000000000101","000000000000010000","111111111111111001","000000000000000000","000000000000000011","111111111111101001","000000000000110000","111111111111100010","000000000000011000","000000000000010000","000000000000010110","000000000000011111","000000000000000111","111111111111110101","000000000000000111","000000000000011010","111111111111011000","111111111111110101","000000000000001000","000000000000001000","000000000000100010","111111111111100101","000000000000000101","111111111111110001","000000000000001111","000000000000001101","111111111111101111","111111111111100001","000000000000000100","111111111111111001","111111111111011001","000000000000001110","111111111111110001","000000000000011111","111111111111011010","111111111111110110","111111111111111110","000000000000101000","000000000000001101","000000000000011000","111111111111111011","000000000000001010","000000000000000000","111111111111101111","111111111111110110","000000000000101000","000000000000001110","000000000000000110","111111111111111101","111111111111010000","111111111111111110","111111111111110110","111111111111101110","000000000000000110","000000000000000001","111111111111100110","000000000000001101","000000000000010101","000000000000100001","000000000000000110","000000000000011111","111111111111110101","000000000000000001","000000000001001111","000000000000000000","000000000000011010","111111111111111011","111111111111100001","000000000000001000","111111111111001011","111111111111100000","000000000000100001","000000000000001111","111111111111111010","000000000000000010","000000000000010000","111111111111110100","111111111111111111","000000000000010110","111111111111111000","000000000000001011","111111111111011110","111111111111100101","000000000000011110","000000000000010110","111111111111111101","111111111111111010","000000000000000100","000000000000011010","111111111111111001","000000000000011100","111111111111100010","000000000000011000","111111111111011001","111111111111100111","000000000000001101","111111111111100111","000000000000011101","000000000000010001","111111111111111100","000000000000110010","000000000000001000","111111111111110011","000000000000010111","000000000000000000","111111111111111100","111111111111101011","000000000000100001","111111111111101011","000000000000100000","000000000000100001","000000000000000010","111111111111100001","000000000000000000","111111111111100010","000000000000001010","000000000000010000","111111111111100110","111111111110010111","000000000000101000","111111111111110101","000000000000011001","111111111111011100"),
("000000000000100001","111111111111011111","000000000000100111","000000000000001001","000000000000001000","000000000000010110","000000000000000110","000000000000001100","111111111111110110","111111111111100000","000000000000000100","000000000000011111","111111111111010111","000000000000011011","111111111111110000","000000000000010001","000000000000010111","000000000000000101","000000000000001000","111111111111101111","000000000000011000","111111111111001101","111111111111101000","111111111111110110","111111111111110101","000000000000001111","000000000000001101","000000000000000010","000000000000000110","000000000000001000","000000000000010011","111111111111110101","111111111111111101","000000000000010100","000000000000010011","111111111111110110","111111111111110010","111111111111100111","000000000000101110","111111111111011001","111111111111100110","000000000000001000","000000000000110011","000000000000010111","000000000000000000","000000000000010011","000000000001000000","111111111111101110","000000000000000001","111111111111101100","000000000000011111","000000000000010011","111111111111101100","111111111111110101","111111111111010111","000000000000001110","111111111111100100","111111111111111010","000000000000000111","111111111111111110","111111111111111000","000000000000000000","000000000000001010","000000000000011111","000000000000010111","111111111111111010","111111111111110101","000000000000100110","000000000000111010","111111111111011000","000000000000011110","111111111111110011","111111111111011000","000000000000000000","111111111111100011","111111111111111000","000000000000011001","111111111111101000","111111111111110110","000000000000010100","000000000000100011","000000000000100001","000000000000000111","000000000000101011","111111111111110110","000000000000001001","111111111111110001","111111111111111000","000000000000101101","000000000000010000","000000000000000011","000000000000010000","000000000000001101","000000000000000011","111111111111111110","000000000000100110","111111111111100000","000000000000001010","000000000000001001","111111111111101100","000000000000101000","000000000000000001","111111111111111001","000000000000001011","000000000000011101","000000000000001111","111111111111110000","000000000000000010","000000000000100100","000000000000010001","000000000000001101","111111111111111100","000000000000101010","111111111111110010","000000000000000100","000000000000000011","000000000000010001","111111111111010111","000000000000000001","111111111111101010","111111111111101110","000000000000101100","000000000000001000","111111111101001011","000000000000101101","000000000000010101","000000000000101010","111111111111110100"),
("000000000000001100","111111111111010100","000000000000011011","111111111111111101","000000000000000001","000000000000001010","000000000000001010","111111111111110111","111111111111110110","111111111111010001","000000000000101101","000000000000011001","000000000000001011","000000000000001001","111111111111101000","000000000000000011","000000000000010100","000000000000011001","000000000000010101","111111111111110100","111111111111111110","000000000000000101","111111111111011111","111111111111111101","111111111111110101","000000000000100100","000000000000011110","000000000000001010","000000000000010010","000000000000000110","111111111111111011","111111111111111000","000000000000010011","111111111111100110","000000000000001010","111111111111111000","111111111111111011","111111111111110011","000000000000101100","000000000000010000","111111111111100011","000000000000100111","000000000000001010","000000000000100000","000000000000010101","111111111111101010","000000000001001111","111111111111110011","111111111111100111","000000000000000000","111111111111010110","000000000000010001","111111111111111111","000000000000001110","111111111111010011","000000000000001000","000000000000001110","111111111111111011","111111111111110001","000000000000000001","111111111111100100","111111111111101101","111111111111111000","000000000000011010","000000000000000000","111111111111101001","111111111111110111","000000000000011101","000000000000111101","111111111111011100","000000000000011001","000000000000000001","111111111111110111","111111111111110111","111111111111010011","111111111111111001","000000000000001000","000000000000001000","111111111111110001","111111111111110101","000000000000000010","000000000000011110","000000000000010100","000000000000010110","111111111111111100","000000000000010101","000000000000001111","111111111111100000","000000000000000001","000000000000010011","111111111111101001","111111111111111111","000000000000011000","000000000000000000","000000000000000101","000000000000001000","111111111110111101","000000000000010010","000000000000000001","111111111111100010","000000000000101000","000000000000001011","111111111111110110","000000000000000000","000000000000011000","000000000000001000","000000000000001001","000000000000001000","000000000000001011","111111111111110110","000000000000010111","000000000000000100","000000000000100001","111111111111110001","000000000000010111","000000000000000000","000000000000011010","111111111111101110","000000000000101100","111111111111110100","000000000000001011","000000000000100010","111111111111110101","111111111101111111","000000000000000000","000000000000001101","000000000000001101","111111111111101110"),
("000000000000001110","111111111111011010","111111111111111110","000000000000010011","000000000000000101","000000000000011111","111111111111110001","000000000000000000","000000000000000001","111111111111010010","000000000000111010","000000000000001100","111111111111111111","000000000000001110","111111111111001110","000000000000000000","000000000000010001","000000000000001101","000000000000011011","000000000000010001","111111111111110011","000000000000001110","111111111111111000","000000000000001011","111111111111111000","000000000000101100","000000000000011100","000000000000010001","000000000000011101","111111111111111101","000000000000010100","111111111111101001","000000000000000101","111111111111111010","000000000000011110","000000000000000101","111111111111111101","000000000000011011","000000000000100000","111111111111101111","111111111111100101","000000000000101010","000000000000000111","000000000000001010","000000000000001101","000000000000000000","000000000000100111","000000000000011011","000000000000001101","000000000000010011","111111111110110011","111111111111111001","111111111111110111","000000000000000011","111111111111101110","000000000000011110","000000000000000111","000000000000001010","111111111111011001","111111111111111001","111111111111011111","000000000000000101","111111111111100101","000000000000001010","111111111111111011","111111111111110111","000000000000001111","000000000000010110","000000000001000001","111111111111101011","000000000000011001","000000000000100000","000000000000001001","000000000000000101","111111111111111000","111111111111101011","000000000000001001","000000000000010001","111111111111110110","000000000000010010","000000000000001101","111111111111110011","000000000000011101","000000000000100001","000000000000001110","111111111111110001","111111111111011111","111111111111101101","000000000000010111","000000000000010001","111111111111101100","111111111111100100","000000000000000001","111111111111111110","111111111111101111","000000000000010001","111111111111011000","000000000000011001","000000000000001100","000000000000010100","000000000000100001","000000000000001011","111111111111110110","111111111111111111","000000000000001101","111111111111111111","000000000000000000","000000000000010000","000000000000100011","111111111111100000","000000000000001100","111111111111111000","000000000000101000","111111111111111111","000000000000100011","000000000000001000","000000000000010011","111111111111100111","000000000000101110","000000000000001100","111111111111110110","000000000000010000","000000000000010011","111111111111010010","000000000000010001","111111111111101100","111111111111111011","000000000000000111"),
("000000000000010011","111111111111101101","000000000000001011","111111111111111100","111111111111110111","000000000000011000","000000000000011101","000000000000001010","000000000000010101","111111111111101110","000000000000100111","000000000000001110","000000000000011101","111111111111111001","111111111111111000","000000000000001100","000000000000001111","000000000000000001","000000000000000110","111111111111110011","111111111111011100","000000000000001010","111111111111010101","000000000000010000","111111111111100110","000000000000011111","111111111111111100","111111111111101001","000000000000101111","000000000000000101","000000000000000000","000000000000010010","111111111111111011","000000000000001010","000000000000010111","111111111111111101","000000000000001010","000000000000011100","000000000000001011","111111111111111100","111111111111100010","000000000000011111","000000000000010011","000000000000010111","000000000000001110","000000000000001010","000000000000110010","000000000000101111","111111111111110010","111111111111110000","111111111111101010","000000000000000000","111111111111101011","000000000000001001","000000000000010000","000000000000011011","000000000000000011","111111111111100101","111111111111111011","111111111111110101","111111111111011011","000000000000000010","111111111111100011","000000000000001101","000000000000000100","111111111111101011","000000000000010101","111111111111110000","000000000000001101","111111111111110011","000000000000100011","000000000000001001","111111111111110001","111111111111110001","000000000000000011","111111111111110111","111111111111111111","000000000000000001","000000000000000111","000000000000010001","000000000000000010","111111111111110010","000000000000010010","000000000000011011","000000000000001111","111111111111110011","111111111111111100","000000000000001000","000000000000010010","000000000000001010","000000000000000111","111111111111100011","111111111111101101","111111111111111011","000000000000001000","111111111111110000","111111111111010001","111111111111110101","111111111111101001","000000000000101000","000000000000010011","000000000000001010","000000000000000110","000000000000000010","000000000000001111","000000000000010111","111111111111111100","000000000000010111","000000000000101011","111111111111110110","111111111111111011","000000000000000000","000000000000001011","000000000000010110","000000000000100101","000000000000000000","000000000000000101","111111111111111101","000000000000010110","111111111111111110","111111111111110001","000000000000000000","000000000000101001","000000000000011110","000000000000011010","000000000000000101","111111111111101110","000000000000000000"),
("000000000000011101","111111111111111010","000000000000010011","000000000000001111","000000000000010111","000000000000001000","000000000000000101","111111111111111011","000000000000000101","111111111111101010","111111111111100011","000000000000000100","000000000000000010","000000000000001000","000000000000010110","111111111111110101","000000000000000000","111111111111110110","111111111111110010","111111111111110000","111111111111101001","111111111111010110","111111111111111011","000000000000000001","000000000000000000","000000000000010101","000000000000010101","111111111111101110","000000000000010101","111111111111110111","000000000000000010","000000000000000001","111111111111110101","111111111111101110","000000000000001001","111111111111110100","000000000000000110","000000000000010111","111111111111111111","000000000000001001","111111111111101110","000000000000001001","000000000000000111","111111111111110010","000000000000001111","000000000000001101","000000000000001011","000000000000110101","000000000000010101","000000000000010100","111111111111111101","000000000000001110","111111111111100001","000000000000000010","000000000000001101","000000000000000100","000000000000000011","111111111111110010","111111111111101010","111111111111101011","111111111111100111","000000000000000100","000000000000000110","111111111111101001","000000000000000111","000000000000010001","000000000000010010","111111111111110110","000000000000010111","111111111111111101","111111111111110010","000000000000001011","000000000000000000","111111111111111000","111111111111101110","111111111111100011","000000000000011010","000000000000001100","000000000000010100","000000000000000010","000000000000001011","111111111111101010","000000000000111000","000000000000010011","111111111111110100","000000000000011100","111111111111110010","111111111111101101","111111111111110101","000000000000000001","000000000000100111","111111111111011001","111111111111111110","111111111111101101","000000000000000110","111111111111110110","111111111111110001","000000000000000101","111111111111100110","111111111111110011","000000000000001011","000000000000011001","000000000000000001","111111111111101101","111111111111011011","000000000000001110","000000000000011001","000000000000101101","000000000000011011","000000000000101100","000000000000000101","111111111111011011","000000000000001111","000000000000010101","000000000000110111","111111111111101101","000000000000000000","111111111111111101","000000000000001101","111111111111111000","111111111111101110","000000000000000001","000000000000100000","000000000001000000","000000000000011100","111111111111110001","111111111111110101","111111111111110001"),
("111111111111111100","111111111110111010","000000000000001100","111111111111110110","000000000000011001","000000000000100111","000000000000000011","111111111111110001","111111111111111111","111111111111011010","111111111111110111","111111111111111101","111111111111111100","000000000000000010","000000000000010000","111111111111111011","000000000000001010","000000000000001010","111111111111111100","000000000000001100","111111111111111001","111111111111011100","111111111111110000","111111111111110010","111111111111110010","000000000000010001","111111111111101100","111111111111110111","111111111111111110","000000000000000000","111111111111111110","111111111111101110","111111111111111111","111111111111111011","000000000000010001","111111111111101100","000000000000000110","111111111111111000","000000000000010101","111111111111100111","111111111111101000","111111111111111010","111111111111110001","000000000000010111","000000000000011010","000000000000000011","000000000000010010","000000000000011000","000000000000010010","111111111111110010","111111111111111010","000000000000000010","111111111111100011","111111111111101110","000000000000010110","000000000000100010","000000000000000000","111111111111101011","111111111111110001","111111111111111011","111111111111110001","111111111111111101","111111111111111110","111111111111110110","000000000000000011","000000000000011001","000000000000010100","111111111111111011","111111111111111000","111111111111110001","000000000000000001","111111111111110011","111111111111111110","000000000000000011","000000000000000110","000000000000010010","000000000000100001","000000000000000101","000000000000001011","000000000000000000","000000000000010010","111111111111110110","000000000001000110","111111111111110010","000000000000000000","000000000000110110","000000000000000000","111111111111110010","000000000000001111","000000000000001100","000000000000010011","111111111111101110","000000000000000110","000000000000000011","000000000000011000","000000000000011101","000000000000100001","111111111111110010","000000000000000101","111111111111101000","000000000000011100","000000000000001100","111111111111110110","000000000000000001","111111111111101001","111111111111110101","000000000000100110","000000000000000111","000000000000100010","000000000000111001","000000000000011111","111111111111011010","000000000000010100","111111111111110010","000000000000100101","000000000000001111","111111111111110010","111111111111101001","000000000000010100","111111111111110010","111111111111110000","111111111111101100","000000000000000100","000000000000010101","000000000000101111","111111111111110101","000000000000001011","000000000000000101"),
("111111111111110111","111111111111010100","000000000000000010","000000000000000101","111111111111110110","111111111111111001","000000000000011100","000000000000000001","111111111111111111","000000000000000000","111111111111100010","111111111111010010","111111111111111100","111111111111110110","000000000000101110","111111111111111011","000000000000011000","111111111111100000","000000000000000110","000000000000010000","111111111111101010","111111111111111011","000000000000000000","111111111111100111","111111111111101100","000000000000001100","111111111111101110","111111111111110100","111111111111101000","111111111111111010","000000000000000001","111111111111100010","000000000000001101","111111111111101101","111111111111100101","111111111111100000","000000000000010001","111111111111111001","000000000000011110","000000000000011010","111111111111111010","111111111111010111","000000000000010000","111111111111111010","000000000000001000","000000000000000000","111111111111101110","000000000000011011","000000000000011111","000000000000010001","000000000000000010","000000000000001011","111111111111110111","000000000000000000","000000000000000100","000000000000010101","000000000000100100","111111111111111010","000000000000011110","000000000000010000","000000000000001001","000000000000010000","000000000000010101","000000000000000000","111111111111011101","000000000000100110","000000000000001111","000000000000000001","111111111111110011","111111111111110110","111111111111110101","111111111111110100","000000000000001001","000000000000010011","111111111111111001","000000000000000011","000000000000010000","111111111111110101","000000000000100001","000000000000010101","000000000000010010","000000000000000100","000000000000101001","000000000000000010","111111111111011111","000000000000101000","000000000000011011","111111111111101001","000000000000010001","111111111111101110","000000000000010100","111111111111100111","000000000000001000","111111111111110100","000000000000110001","000000000000000101","000000000000000100","000000000000101110","000000000000001000","111111111111111011","000000000000011101","111111111111111001","000000000000000111","111111111111110111","111111111111110000","000000000000010010","000000000000011001","000000000000010001","000000000000000111","000000000000101110","000000000000010101","111111111111011010","000000000000000000","000000000000010110","111111111111111110","000000000000000011","000000000000000000","111111111111110111","000000000000001011","111111111111101110","111111111111101010","000000000000000000","111111111111101101","000000000000000001","000000000000110100","000000000000000100","111111111111110111","000000000000010100"),
("111111111111100101","111111111111111100","000000000000000010","111111111111101000","000000000000001011","000000000000000100","000000000000000101","000000000000010011","111111111111100111","000000000000001010","111111111111100111","111111111111011111","000000000000000010","111111111111101111","000000000000101010","111111111111011110","000000000000100000","111111111111010110","111111111111111101","000000000000001010","000000000000000011","111111111111110100","000000000000000111","111111111111100111","111111111111101111","111111111111110011","111111111111101111","111111111111101100","000000000000011001","000000000000001001","111111111111110000","000000000000001100","000000000000000000","000000000000010000","111111111111100111","111111111111101010","111111111111110100","000000000000000100","000000000000001010","000000000000100101","111111111111110011","111111111111111101","111111111111110010","000000000000000001","000000000000011000","000000000000001011","000000000000000010","000000000000000000","000000000000010011","000000000000000000","000000000000001001","111111111111111110","111111111111100110","000000000000011001","111111111111110100","000000000000010111","000000000000001011","000000000000001100","111111111111111111","111111111111110011","000000000000010010","000000000000001000","111111111111110011","000000000000001111","111111111111000010","000000000000011111","111111111111101101","111111111111111111","000000000000011000","111111111111101010","111111111111111001","000000000000000110","000000000000001100","000000000000010101","000000000000011100","111111111111111111","000000000000010000","000000000000000101","000000000000100000","000000000000011010","111111111111111111","000000000000000100","000000000000110001","000000000000001110","111111111111110011","000000000000111001","000000000000001101","111111111111111110","111111111111111001","000000000000010000","000000000000001110","000000000000000001","111111111111101011","000000000000001111","000000000000001010","111111111111111011","000000000000010111","000000000000100100","000000000000011000","111111111111111101","111111111111110000","111111111111110011","111111111111110101","111111111111100000","000000000000000010","111111111111101110","111111111111110100","000000000000001001","000000000000001001","000000000000010110","111111111111111101","111111111111111011","000000000000010101","000000000000001010","111111111111111100","111111111111110101","111111111111111011","111111111111111101","000000000000001000","111111111111110100","111111111111111100","111111111111110100","111111111111010111","111111111111100100","000000000000001110","111111111111101111","111111111111100010","000000000000001011"),
("111111111111101000","111111111111101100","000000000000000001","111111111111100111","000000000000011100","111111111111101001","000000000000010101","111111111111111001","111111111111101011","000000000000000000","111111111111100111","111111111111101001","000000000000000001","111111111111110101","000000000000011110","111111111111110010","000000000000011000","111111111111110010","000000000000010100","000000000000000001","111111111111101101","000000000000000101","111111111111111100","111111111111100000","000000000000001010","111111111111111001","000000000000001000","111111111111011010","000000000000001111","111111111111111000","111111111111110000","000000000000000001","000000000000001101","111111111111111101","111111111111011011","111111111111100011","000000000000010110","000000000000001001","111111111111111101","000000000000100110","111111111111110110","000000000000000000","000000000000010100","111111111111110111","000000000000001100","111111111111110100","000000000000010000","000000000000000010","000000000000100100","111111111111110000","000000000000010100","111111111111101101","111111111111110100","000000000000001100","111111111111111100","111111111111110110","000000000000000111","000000000000000111","000000000000001000","000000000000010010","111111111111111010","111111111111111000","111111111111110111","000000000000000001","111111111110101010","111111111111111011","111111111111010011","000000000000001100","000000000000011001","111111111111110100","111111111111110101","000000000000010010","111111111111111111","000000000000010000","000000000000011001","000000000000100001","111111111111111001","111111111111100010","000000000000101001","000000000000000001","111111111111100001","111111111111111010","000000000000010100","000000000000101110","111111111111111101","000000000000110001","000000000000010111","000000000000000000","000000000000000010","000000000000001101","000000000000001000","111111111111111111","000000000000000010","000000000000010011","111111111111110100","111111111111111001","000000000000010100","000000000000101011","000000000000011110","000000000000000000","000000000000000101","111111111111111000","111111111111110101","111111111111110001","111111111111110110","111111111111101110","111111111111011111","111111111111110101","111111111111101010","000000000000000111","111111111111101111","000000000000100001","000000000000000101","000000000000011110","111111111111110111","000000000000000000","000000000000011000","000000000000001110","111111111111101010","000000000000000000","000000000000001110","000000000000000100","111111111111010000","111111111111110011","000000000000010011","111111111111111101","111111111111010101","111111111111110001"),
("111111111111100110","000000000000001110","000000000000010001","111111111111000111","000000000000001010","000000000000000010","000000000000001101","000000000000010010","111111111111110110","000000000000000111","111111111111010000","000000000000001001","000000000000000001","111111111111101100","000000000000011000","111111111111111111","000000000000000010","111111111111101010","000000000000000000","111111111111101111","111111111111101010","000000000000010111","111111111111111101","111111111111111000","111111111111111010","111111111111101101","111111111111100011","111111111111111111","000000000000011010","111111111111101011","000000000000001100","111111111111111011","000000000000001110","000000000000001100","111111111111110001","111111111111110100","000000000000011001","000000000000001011","111111111111101001","000000000000101000","000000000000000100","000000000000000010","000000000000001100","111111111111010100","000000000000010101","000000000000000111","111111111111111101","111111111111110111","000000000000100100","111111111111110000","000000000000001001","111111111111111001","111111111111110101","000000000000010001","000000000000001010","111111111111110100","111111111111101101","000000000000001101","000000000000010000","111111111111110011","000000000000011001","000000000000000001","111111111111111100","111111111111110011","111111111111110011","111111111111111111","111111111111100101","000000000000000000","000000000000000000","111111111111011011","111111111111111000","000000000000000110","000000000000000110","000000000000001110","111111111111111111","000000000000010101","000000000000000000","111111111111110010","000000000000011000","000000000000010111","111111111111100110","000000000000010011","000000000000101111","111111111111111101","111111111111101110","111111111111111101","000000000000000111","000000000000011011","111111111111101101","000000000000001100","000000000000000110","111111111111111000","111111111111101001","000000000000000011","111111111111111101","111111111111011101","000000000000010111","000000000000010101","000000000000011010","111111111111111101","111111111111110001","111111111111101000","111111111111101001","111111111111110110","111111111111011111","111111111111100101","111111111111101000","000000000000000110","111111111111011001","000000000000100001","111111111111101100","000000000000001110","111111111111110011","000000000000000111","111111111111101101","111111111111111011","111111111111110111","111111111111111101","111111111111100011","000000000000010100","000000000000001011","111111111111101011","111111111111110000","111111111111110110","000000000000000000","000000000000010010","111111111111100101","000000000000001000"),
("111111111111111011","111111111111111110","111111111111111001","111111111111100110","000000000000000110","000000000000001110","000000000000000001","000000000000000101","111111111111101010","111111111111111000","111111111111111011","000000000000000000","000000000000001100","111111111111101000","111111111111111111","000000000000011100","000000000000010000","111111111111110101","111111111111111001","000000000000011011","000000000000000010","000000000000101001","000000000000000100","111111111111111100","000000000000001100","111111111111111100","111111111111100110","111111111111101111","000000000000010100","111111111111000101","111111111111110100","111111111111110010","000000000000001000","111111111111111010","111111111111111010","111111111111111000","000000000000001111","000000000000000101","111111111111100111","000000000000001000","000000000000010001","000000000000010101","111111111111111100","111111111111101111","000000000000001100","000000000000010111","000000000000001100","000000000000010100","000000000000000010","111111111111101010","000000000000011011","111111111111111111","000000000000001100","000000000000000110","000000000000001000","000000000000000000","111111111111010001","111111111111101111","000000000000000111","111111111111110101","111111111111110011","000000000000000001","000000000000010000","111111111111111101","000000000000010000","000000000000001010","111111111111000101","111111111111110011","000000000000011110","111111111111110101","111111111111111011","111111111111100110","111111111111001110","000000000000010010","000000000000010010","000000000000111101","000000000000010111","000000000000000101","000000000000000110","000000000000011000","111111111111110110","111111111111100000","000000000001000101","111111111111011110","111111111111101011","111111111111111011","111111111111111010","000000000000110111","111111111111110101","000000000000001110","000000000000000001","111111111111011110","111111111111111001","000000000000010011","111111111111110110","111111111111000100","000000000000000010","000000000000001110","000000000000001001","111111111111100010","000000000000100100","111111111111011000","111111111111011111","111111111111100011","111111111111111100","111111111111111010","111111111111111001","111111111111110000","111111111111110101","111111111111111100","111111111111111110","111111111111111010","111111111111110100","111111111111111011","000000000000000000","111111111111101010","111111111111111001","000000000000011000","111111111111000110","000000000000000101","000000000000010011","000000000000000010","111111111111111010","000000000000011001","000000000000100010","000000000000001101","111111111111110000","111111111111011010"),
("000000000000000111","000000000000101011","111111111111111100","111111111111011100","111111111111101001","111111111111110101","111111111111110100","111111111111111110","000000000000010001","000000000000001011","111111111111111000","000000000000011100","111111111111101010","111111111111110011","111111111111111010","000000000000011010","111111111111110011","111111111111110110","111111111111101011","000000000000000010","111111111111111000","000000000000001010","111111111111110010","111111111111101011","111111111111101111","111111111111111111","000000000000000110","000000000000000111","000000000000001010","111111111111011100","111111111111100111","000000000000001010","111111111111111101","111111111111101000","111111111111100110","111111111111110101","000000000000011111","000000000000001010","111111111111010001","000000000000010101","000000000000000100","000000000000010000","000000000000000000","111111111111101100","000000000000000010","000000000000010000","000000000000001101","111111111111110100","111111111111111100","111111111111111111","111111111111111101","111111111111111000","111111111111111011","000000000000010000","000000000000001101","000000000000001001","111111111111100001","000000000000001010","111111111111101001","000000000000001101","000000000000000001","111111111111110101","111111111111101010","111111111111110100","000000000000001100","111111111111111101","111111111110111000","000000000000000000","000000000000101111","000000000000000000","000000000000001111","111111111111111110","111111111111011101","000000000000011101","111111111111111001","000000000001000010","000000000000001011","000000000000001010","000000000000000101","000000000000011100","111111111111101010","000000000000000001","000000000000010011","111111111111000011","000000000000001010","111111111111110010","000000000000001111","000000000000100010","000000000000001010","000000000000010010","111111111111101010","000000000000011000","000000000000001000","000000000000001010","111111111111101100","000000000000000000","000000000000010011","000000000000100000","111111111111110001","000000000000001100","111111111111111011","111111111111111100","000000000000010000","111111111111011111","111111111111101111","000000000000000100","111111111111110110","000000000000010010","111111111111101001","000000000000001010","111111111111111101","111111111111101100","111111111111111111","000000000000011011","111111111111111010","000000000000001010","000000000000000110","000000000000000011","111111111111011001","000000000000010111","111111111111111111","000000000000000011","000000000000000011","000000000000000000","000000000000100101","111111111111110111","000000000000001101","111111111111110001"),
("111111111111101110","000000000000100000","000000000000000101","111111111111111100","000000000000000000","000000000000001001","111111111111101111","000000000000000111","111111111111111110","111111111111111101","000000000000000001","000000000000011010","111111111111111100","111111111111010100","111111111111101000","000000000000010111","111111111111111000","111111111111101101","111111111111100010","000000000000000001","000000000000000011","000000000000001001","111111111111111011","111111111111110000","111111111111111101","111111111111111000","111111111111111100","000000000000001010","000000000000001110","111111111111110100","111111111111110100","111111111111101010","000000000000000110","111111111111010010","111111111111101111","111111111111111111","111111111111101101","000000000000010000","111111111110110111","111111111111111110","111111111111111010","111111111111111010","000000000000001000","111111111111100110","000000000000001101","111111111111110011","000000000000010110","000000000000010111","000000000000000101","111111111111110011","000000000000010100","111111111111110101","000000000000010101","111111111111101000","000000000000001101","111111111111110000","111111111111011001","111111111111101101","111111111111101101","111111111111110010","111111111111101101","111111111111001010","000000000000001110","111111111111100010","000000000000001001","111111111111111111","111111111110101010","000000000000010010","000000000000110101","000000000000000001","111111111111111010","111111111111110000","111111111110111110","000000000000010001","000000000000001000","000000000000110000","000000000000001110","111111111111110111","111111111111101001","000000000000010101","111111111111101010","111111111111011100","000000000000001111","111111111110111101","000000000000001100","111111111111110011","000000000000001100","000000000000010011","111111111111101111","000000000000010000","000000000000000001","000000000000010001","000000000000001000","000000000000000101","000000000000001010","111111111111101001","000000000000110110","000000000000011011","111111111110111000","111111111111101010","111111111111111100","111111111111110110","111111111111100101","111111111111111001","111111111111111011","000000000000011100","111111111111110100","111111111111101110","111111111111010110","111111111111100100","000000000000010010","111111111111000100","000000000000001100","000000000000100011","111111111111111100","111111111111111010","000000000000001111","111111111111110001","111111111111000111","111111111111111111","111111111111101010","000000000000001110","000000000000000000","000000000000001000","000000000000010011","000000000000000111","000000000000001100","000000000000000110"),
("111111111111110000","000000000000011100","111111111111111101","111111111111100111","000000000000000000","111111111111111110","111111111111100011","000000000000011101","000000000000000101","000000000000011001","000000000000100111","000000000000101101","111111111111111111","111111111111010010","111111111111011010","000000000000110111","000000000000001000","111111111111111110","111111111111011010","000000000000011111","000000000000010000","000000000000011010","111111111111111100","000000000000000111","111111111111111011","000000000000011000","111111111111101000","111111111111111100","000000000000011110","111111111111101111","000000000000000000","111111111111111011","111111111111111101","111111111111010111","111111111111100000","000000000000000100","000000000000001111","000000000000010111","111111111110111001","000000000000011111","000000000000011101","111111111111110000","000000000000011000","111111111111110010","111111111111111111","111111111111100000","000000000000010111","000000000000000000","000000000000000100","000000000000000000","000000000000100000","111111111111111011","111111111111110100","000000000000000000","000000000000010111","111111111111101011","111111111111001010","111111111111111111","111111111111111011","000000000000000101","111111111111100101","111111111111111101","111111111111111100","111111111111100001","000000000000001001","111111111111011000","111111111111101001","000000000000010000","000000000000011101","111111111111111110","000000000000001001","111111111111111010","111111111110110100","000000000000001001","000000000000001010","000000000000101010","111111111111110010","111111111111111011","111111111111010110","000000000000000100","111111111111110000","111111111111011101","000000000000011101","111111111111001000","000000000000000000","111111111111001001","000000000000001110","000000000000011011","111111111111111011","000000000000011110","111111111111110110","111111111111111100","000000000000000110","111111111111111011","000000000000000011","111111111111110010","000000000000010010","111111111111101100","111111111111101010","111111111111110000","111111111111100001","111111111111111001","111111111111100010","000000000000001000","000000000000010100","000000000000101101","111111111111101110","000000000000000101","111111111111011101","111111111111110100","111111111111011001","111111111111101111","000000000000010011","000000000000010001","111111111111110000","000000000000001000","000000000000000001","000000000000001111","111111111111100101","000000000000000110","111111111111110000","111111111111111010","000000000000001100","111111111111110111","000000000000011001","111111111111110000","000000000000001110","111111111111111100"),
("000000000000110001","000000000000011010","111111111111101010","000000000000001000","000000000000010011","000000000001010110","000000000000110001","000000000000000001","111111111111101111","111111111111101100","000000000000101111","000000000000000101","111111111111110011","111111111111000000","111111111111101111","000000000000100010","000000000000000011","111111111111111000","111111111111101011","000000000000100001","000000000000000011","111111111111111111","111111111111110111","111111111111011011","111111111111010101","000000000000111011","111111111111111000","000000000000001010","111111111111110011","111111111111111000","000000000000011110","111111111111111001","000000000000000000","111111111111101010","000000000000011101","111111111111110001","111111111111111010","000000000000010010","111111111111001101","111111111111100001","111111111111011100","111111111111110100","000000000000111000","000000000000101010","000000000000000000","111111111111010011","000000000000011100","000000000001010000","111111111111001010","111111111111101111","111111111111110101","111111111111111010","111111111111011000","111111111111011101","000000000000000001","111111111111111110","111111111111011110","111111111111101000","111111111110111001","000000000000000000","111111111111010111","111111111111010110","000000000000001000","111111111111110101","111111111111010110","111111111111010010","000000000000001000","000000000000100001","000000000000000101","111111111111100011","000000000000111001","111111111111101010","111111111111101001","111111111111101000","111111111111111110","000000000000111001","000000000001000001","000000000000000000","111111111111100000","000000000000011101","111111111111100101","000000000000010000","000000000000110001","111111111111011010","111111111111100001","111111111111100111","000000000000001000","000000000000010010","111111111111101101","111111111110111001","111111111111111110","111111111111100000","000000000000010100","000000000000101011","111111111111101101","111111111111110111","000000000000000110","000000000000010100","111111111111010011","111111111111100010","000000000001000100","000000000000000000","111111111111001110","111111111111110000","111111111111111111","000000000000100011","111111111111010001","000000000000001111","111111111111001100","111111111111110111","111111111111000010","111111111111110000","000000000000101001","111111111111000011","111111111111000111","000000000000000110","000000000000000100","111111111111110111","111111111111001011","111111111111011010","000000000000110001","000000000001011011","000000000000001100","000000000000000100","000000000000100100","000000000000001001","000000000000011111","111111111111100101"),
("000000000000101011","111111111111100110","000000000000000001","000000000000000111","000000000000000110","000000000001000011","000000000000101011","000000000000101011","000000000000001011","111111111111000110","000000000000100001","111111111111001000","000000000000001000","111111111111110010","111111111111010100","000000000000001101","000000000000001100","000000000000010010","111111111111011100","000000000000100011","000000000000001101","111111111111111111","000000000000000100","111111111111100011","111111111111000001","000000000000100011","111111111111111010","000000000000011001","000000000000010100","111111111111100110","000000000000011010","111111111111101111","000000000000000010","111111111111010000","000000000000111101","000000000000001001","000000000000110110","000000000000110100","111111111111010101","111111111111011010","111111111111010111","111111111111100011","000000000000001000","000000000000011101","000000000000000000","111111111111000000","111111111111101101","000000000000110101","111111111111011110","111111111111100111","111111111111101111","000000000000111001","111111111111011001","111111111111111001","000000000000110110","000000000000100000","111111111111011111","000000000000000000","111111111111000100","000000000000000000","111111111111001110","000000000000010010","000000000000100010","111111111111101101","000000000000000010","111111111111001000","111111111111110111","111111111111101110","000000000000101100","111111111111101001","000000000000000100","000000000000010011","111111111111110101","000000000000010001","111111111111100011","000000000000010101","000000000000100011","000000000000000000","111111111111110011","000000000000110010","111111111111101010","111111111111111010","000000000001001000","000000000000001100","111111111111111110","111111111111011111","000000000000001111","000000000000000010","111111111110111110","111111111111010011","111111111110110100","111111111111010111","111111111111010110","000000000000100000","111111111111111001","111111111111011111","111111111111100000","000000000000001010","111111111111011001","000000000000001101","000000000000101101","111111111111011000","111111111111101000","111111111111111000","000000000000001100","000000000000011101","000000000000000000","111111111111010000","111111111111100111","111111111111011101","111111111111111001","000000000000010100","111111111111101011","111111111111011001","111111111111111111","000000000000101001","111111111111010111","000000000000010000","111111111111001110","111111111111111001","000000000000000110","000000000001011110","000000000000000110","000000000000001111","000000000000110010","111111111111011110","000000000000010100","000000000000001111"),
("000000000000001101","111111111111011001","111111111111100111","000000000000000101","111111111111100011","000000000000000110","000000000000010110","000000000000100101","000000000000011001","111111111111110000","000000000000010011","111111111111010101","000000000000100100","111111111111110111","111111111111011101","000000000000100101","000000000000010101","000000000000000000","111111111111100101","000000000000000101","000000000000000111","000000000000001000","111111111111111000","111111111111110101","111111111111110111","000000000000011111","111111111111110100","000000000000001000","111111111111110011","111111111111101000","000000000000010100","111111111111110110","000000000000100101","111111111111111000","000000000000001001","111111111111101000","000000000000011010","000000000000010010","111111111111100011","111111111111011010","111111111111111100","111111111111110000","000000000000011001","000000000000100110","000000000000000100","111111111111100001","111111111111101011","111111111111110110","111111111111011011","111111111111010111","000000000000001001","000000000000010010","111111111111101000","000000000000000101","000000000000100011","111111111111111110","111111111111110001","000000000000100100","111111111111111010","111111111111111111","111111111111110110","000000000000001110","000000000000011000","111111111111101010","111111111111100011","111111111111110000","000000000000010010","111111111111110000","000000000000001111","111111111111100111","000000000000101100","000000000000011000","000000000000000000","000000000000101000","111111111111011111","000000000000001101","000000000000011000","000000000000001111","111111111111000011","000000000000000000","111111111111101100","000000000000000111","000000000000010111","111111111111010000","000000000000000000","111111111111100011","000000000000001111","111111111111101111","111111111111110000","111111111111100101","111111111111010100","111111111111100011","111111111111011011","000000000000101111","111111111111111110","000000000000000110","000000000000100110","000000000000000001","111111111111011100","111111111111111110","000000000000010101","111111111111100001","111111111111110101","111111111111111011","000000000000000111","000000000000011111","111111111111101100","000000000000000000","111111111111100010","000000000000000000","111111111111110010","000000000000010111","111111111111010110","000000000000000010","111111111111101010","000000000000011101","111111111111111011","000000000000100111","111111111111111011","000000000000011111","000000000000101000","000000000000010100","000000000000101111","000000000000010010","000000000000010101","111111111111110001","000000000000100100","111111111111011001"),
("111111111111111001","111111111111110100","000000000000000111","000000000000000101","000000000000000010","000000000000000111","000000000000000010","000000000000000111","111111111111101111","000000000000001110","000000000000001010","111111111111110110","000000000000010010","111111111111111011","000000000000000011","000000000000000100","000000000000001011","000000000000000111","111111111111110110","000000000000001101","000000000000010001","000000000000001010","111111111111101110","000000000000001000","000000000000010011","000000000000001111","000000000000000000","000000000000010001","000000000000001111","111111111111110111","111111111111110101","111111111111110010","111111111111101111","111111111111101111","111111111111110100","000000000000010001","111111111111111110","000000000000001101","000000000000000111","111111111111111010","111111111111101110","111111111111111001","000000000000010010","111111111111110110","000000000000001100","000000000000000000","000000000000010011","000000000000000110","111111111111110110","111111111111101110","111111111111110000","000000000000001011","111111111111111101","111111111111111000","000000000000010010","111111111111111111","000000000000000110","111111111111111000","111111111111110101","111111111111111110","111111111111111000","000000000000000001","000000000000001110","000000000000001000","000000000000001111","111111111111111001","111111111111110010","000000000000000010","000000000000001111","111111111111111011","000000000000010010","000000000000001010","000000000000001000","000000000000000111","111111111111110001","111111111111110101","111111111111101100","111111111111110001","111111111111101101","000000000000010011","111111111111111110","000000000000001010","111111111111110011","111111111111111110","000000000000001000","000000000000000011","000000000000000011","000000000000001110","000000000000000111","111111111111111110","111111111111101101","000000000000001111","111111111111111101","000000000000000110","000000000000001111","111111111111110111","111111111111110100","000000000000001101","000000000000001000","111111111111110110","111111111111111010","111111111111110000","000000000000000110","000000000000010010","111111111111110010","111111111111111000","000000000000000000","000000000000001110","111111111111111011","111111111111110100","111111111111110011","111111111111111000","000000000000010011","111111111111110000","111111111111110011","000000000000000100","000000000000001100","000000000000001000","000000000000000101","111111111111110000","000000000000010001","000000000000000111","000000000000001001","111111111111110101","000000000000001110","111111111111110000","000000000000010001","111111111111111001"),
("111111111111100101","111111111111111000","111111111111111111","111111111111110001","000000000000010101","000000000000000100","111111111111101011","000000000000000110","000000000000001101","111111111111110110","000000000000000111","000000000000000111","000000000000001010","111111111111111111","111111111111101000","000000000000000001","000000000000001000","000000000000000000","000000000000010110","000000000000000111","111111111111110111","111111111111101111","000000000000000001","111111111111100101","111111111111100010","000000000000000000","111111111111101110","000000000000000110","000000000000000101","000000000000100000","111111111111111011","000000000000100000","111111111111111011","111111111111110001","000000000000000101","000000000000001111","111111111111100000","000000000000100001","000000000000011010","000000000000011001","000000000000000010","111111111111110111","000000000000010010","111111111111110101","111111111111110010","111111111111110011","111111111111110101","111111111111011110","111111111111111011","000000000000010000","111111111111111100","000000000000000100","111111111111100111","000000000000001110","000000000000010011","111111111111110100","000000000000001010","000000000000001001","000000000000000111","111111111111111010","000000000000010100","000000000000001101","000000000000000010","000000000000001100","000000000000011100","111111111111111010","111111111111101110","000000000000001111","000000000000001010","111111111111101100","000000000000001110","000000000000001000","000000000000010110","000000000000010011","000000000000001011","111111111111111000","111111111111100010","111111111111111110","111111111111111111","111111111111101101","111111111111101101","111111111111111101","000000000000001000","000000000000010000","111111111111111110","111111111111101101","111111111111101010","000000000000011001","111111111111111001","000000000000010100","111111111111100110","111111111111110110","000000000000010010","111111111111110000","111111111111011100","000000000000011110","111111111111111011","111111111111111000","000000000000000110","000000000000100000","111111111111101110","000000000000000010","000000000000010001","000000000000000010","111111111111110100","111111111111100011","000000000000010111","000000000000000011","000000000000001110","111111111111110001","111111111111101001","111111111111110100","000000000000000100","000000000000001000","000000000000011110","000000000000011001","000000000000000110","000000000000100001","000000000000010111","000000000000100000","111111111111110010","000000000000000111","000000000000000101","111111111111111001","000000000000001010","111111111111101111","111111111111100010","000000000000001000"),
("000000000000000010","000000000000001100","000000000000001111","000000000000001001","000000000000001111","000000000000011000","111111111111111010","000000000000001011","000000000000001111","000000000000000101","111111111111011100","000000000000100011","111111111111111101","111111111111100111","000000000000000101","111111111111110111","000000000000101010","000000000000001000","000000000000001001","000000000000010110","111111111111001010","111111111111111001","000000000000000111","111111111111111110","111111111111011010","000000000000000111","000000000000000100","111111111111111000","000000000000100101","000000000000000101","111111111111101110","111111111111111101","000000000000001001","111111111111010001","000000000000000011","000000000000001110","111111111111110111","000000000000011011","111111111111101010","000000000000010111","111111111111101001","111111111111011000","111111111111111000","111111111111111100","000000000000001010","111111111111101101","000000000000011011","000000000000011010","111111111111101110","000000000000011011","111111111111110111","000000000000011011","111111111111010110","000000000000000001","000000000000000000","000000000000100101","111111111111111101","000000000000001110","111111111111101110","111111111111110101","000000000000000001","000000000000011001","000000000000011100","000000000000000111","000000000000001011","111111111111011000","111111111111011001","111111111111110011","000000000000000110","000000000000000000","000000000000001000","000000000000001100","111111111111101101","111111111111101010","000000000000000011","000000000000011100","111111111111111001","111111111111101000","111111111111111111","000000000000111100","111111111111110000","111111111111111110","000000000000010001","000000000000000011","000000000000000000","000000000000001100","000000000000011100","000000000000000001","000000000000011101","000000000000001001","000000000000010011","111111111111110010","111111111111110111","000000000000001000","111111111111101001","111111111111101000","000000000000000100","111111111111111101","000000000000000111","111111111111110010","111111111111111011","111111111111110001","111111111111111111","000000000000000010","111111111111101110","000000000000001111","111111111111110110","111111111111100100","111111111111111101","111111111111111100","111111111111111010","000000000000000001","000000000000011111","000000000000001111","000000000000101000","111111111111111000","000000000000000011","000000000000001010","111111111111111100","000000000000001000","111111111111100011","111111111111101111","111111111111111000","000000000000011001","000000000000101100","111111111111100000","111111111111110101","000000000000001001"),
("000000000000011101","000000000000000110","111111111111101000","000000000000000110","111111111111111100","000000000000001010","111111111111110110","111111111111111111","000000000000010000","111111111111101110","111111111111001110","000000000000000001","000000000000000110","111111111111001101","111111111111011100","111111111111101001","000000000000100011","000000000000000010","000000000000011100","000000000000101011","111111111111100100","111111111111100101","111111111111010010","111111111111101100","111111111111101010","000000000000100010","111111111111110011","000000000000001011","000000000000000100","000000000000011011","000000000000110001","000000000000011001","000000000000100100","000000000000011000","000000000000001101","111111111111011001","111111111111110101","000000000000111110","111111111111010100","000000000000011010","000000000000000101","000000000000000001","111111111111110111","111111111111111011","000000000000100100","111111111111101011","111111111111111100","000000000000001101","111111111111111101","111111111111111010","000000000000010011","000000000000111001","111111111111100111","111111111111110011","000000000000010010","000000000000001101","111111111111011101","000000000000001010","111111111111011010","000000000000001000","000000000000001001","000000000000101101","000000000000011000","111111111111101101","111111111111110111","111111111111100110","000000000000000011","000000000000001011","111111111111100010","111111111111111001","000000000000010110","000000000000101011","111111111111110010","111111111111110001","000000000000100111","111111111111101001","000000000000000010","000000000000001000","111111111111101000","000000000000000000","111111111111101101","000000000000101100","000000000000000101","111111111111110010","000000000000011100","111111111111100000","000000000000000100","000000000000010011","111111111111101000","000000000000000100","111111111111111101","000000000000000010","111111111111110111","111111111111110100","111111111111010101","000000000000000011","000000000000010111","000000000000101100","000000000000010011","111111111111110010","000000000000000111","111111111111110110","000000000000000101","000000000000011111","111111111111100111","000000000000000110","111111111111101111","111111111111100001","111111111111111101","111111111111010111","111111111111011100","111111111111111010","000000000000100100","000000000000000101","000000000000111100","111111111111111110","000000000000011000","000000000000100010","000000000000000000","000000000000011001","000000000000001001","111111111111111000","000000000000000010","111111111111110110","000000000000010011","111111111111101101","111111111111111001","000000000000001100"),
("000000000000001101","111111111111111011","111111111111010110","111111111111111111","000000000000011001","000000000000001000","111111111111111100","000000000000001001","111111111111101001","000000000000001011","111111111110111000","111111111111010100","111111111111111001","111111111111011110","000000000000010010","000000000000001111","000000000000100010","000000000000000111","111111111111110001","000000000000100000","111111111111110111","000000000000011011","000000000000001111","111111111111101100","111111111111101111","000000000000010001","000000000000000001","000000000000001100","000000000000001111","000000000000010010","000000000000000111","111111111111110000","000000000000011010","111111111111111101","111111111111110100","111111111111100100","000000000000001010","000000000000011000","111111111111100010","000000000000001000","111111111111101110","111111111111110011","000000000000000000","111111111111110110","111111111111110111","111111111111110000","000000000000010001","000000000000011011","111111111111111011","000000000000000000","000000000000101110","000000000000100111","000000000000001010","111111111111100111","111111111111101110","111111111111111100","000000000000000000","000000000000000011","000000000000010100","111111111111110010","000000000000000000","000000000000101100","000000000000000110","111111111111100101","000000000000000010","111111111111100001","111111111111111101","111111111111111001","111111111111001101","111111111111111011","000000000000000011","000000000000001101","000000000000010101","111111111111110101","000000000000000010","111111111111011001","000000000000010011","111111111111111011","111111111111101010","000000000000011001","111111111111101101","000000000000001011","000000000000010110","111111111111110110","000000000000011111","111111111111101000","111111111111010110","000000000000010100","111111111111110110","000000000000000000","111111111111110101","111111111111111100","000000000000000100","000000000000001111","111111111111011011","111111111111110100","111111111111111100","000000000000010100","000000000000110001","000000000000010000","111111111111110010","111111111111010111","111111111111101110","111111111111111001","111111111111100010","111111111111111111","111111111111010001","111111111111101000","111111111111101011","000000000000000010","111111111111010111","000000000000000100","111111111111111011","000000000000000100","000000000000010111","111111111111101100","111111111111101111","111111111111110011","111111111111101110","111111111111111101","111111111111101011","111111111111011001","111111111111111110","111111111111110101","000000000000010111","111111111111110010","111111111111111000","111111111111110000"),
("000000000000000110","000000000000010100","111111111111110101","000000000000000011","111111111111111110","111111111111111001","111111111111101101","111111111111110011","111111111111100011","111111111111110011","111111111110101111","111111111111110011","111111111111011001","000000000000010100","000000000000000010","000000000000010101","000000000000001111","111111111111111001","111111111111011101","000000000000010000","000000000000010111","000000000000010110","000000000000010010","111111111111100000","000000000000100000","111111111111110110","111111111111110000","111111111111111000","111111111111111010","111111111111100001","000000000000100110","000000000000001011","000000000000000000","000000000000000010","111111111111111001","111111111111011000","000000000000000011","000000000000001101","111111111111011011","111111111111111110","111111111111011111","111111111111011000","000000000000001011","111111111111000011","111111111111110111","111111111111110001","111111111111111101","000000000000000110","111111111111110011","111111111111111011","000000000000010001","000000000000010001","000000000000000010","111111111111010001","111111111111101111","000000000000000100","111111111111101101","000000000000001110","111111111111111001","111111111111101011","000000000000000011","000000000000010101","111111111111110100","111111111111011111","000000000000010000","111111111111110011","000000000000110000","111111111111101110","000000000000010000","000000000000011001","111111111111111011","111111111111111111","000000000000101100","111111111111011100","000000000000000100","111111111111000101","000000000000011110","111111111111111001","000000000000000001","000000000000001101","111111111111110000","000000000000011001","000000000000011100","111111111111110111","111111111111110000","111111111111110100","111111111111010000","000000000000010110","111111111111100101","111111111111110000","111111111111110101","111111111111101001","000000000000001001","000000000000001001","111111111111010110","111111111111110100","111111111111100110","000000000000001000","000000000000010011","000000000000001001","111111111111110010","111111111111100010","111111111111110111","111111111111111000","000000000000001101","000000000000001111","111111111111000111","111111111111110011","111111111111010111","000000000000000111","111111111111011111","111111111111111111","111111111111111100","000000000000010010","000000000000100010","111111111111111010","111111111111110011","111111111111011110","111111111111010100","111111111111011110","111111111111101111","111111111111101111","111111111111101011","111111111111100000","000000000000010000","111111111111110100","000000000000001011","111111111111101011"),
("000000000000011111","000000000000101111","000000000000001101","000000000000001000","111111111111111100","000000000000011011","000000000000000111","111111111111101101","111111111111111111","000000000000000010","111111111110100000","111111111111101110","111111111111111100","111111111111101101","000000000000001101","000000000000001111","000000000000000001","000000000000010001","111111111111011101","000000000000001010","000000000000010111","000000000000100010","000000000000001111","111111111111110101","000000000000010011","000000000000011011","111111111111100101","111111111111111111","000000000000010100","111111111111000111","000000000000011010","111111111111110010","000000000000011011","111111111111110110","111111111111100001","111111111111100011","000000000000000111","000000000000011100","111111111111011111","111111111111111110","111111111111010110","000000000000001000","111111111111111011","111111111110110110","111111111111111100","111111111111110110","111111111111101101","000000000000010111","111111111111110001","111111111111011001","000000000000000011","000000000000000110","000000000000010010","111111111111100010","111111111111100011","000000000000100011","111111111111101001","111111111111111011","111111111111111101","111111111111110000","000000000000000100","000000000000010110","000000000000001100","111111111111101010","111111111111000011","000000000000000100","000000000000100000","111111111111100000","000000000000000101","000000000000010000","111111111111111011","111111111111100100","000000000000011111","111111111111101010","000000000000001011","111111111111101001","000000000000100001","111111111111110001","000000000000001000","111111111111111101","111111111111101101","000000000000001010","000000000000100000","111111111111011111","111111111111111001","111111111111100110","111111111110101001","111111111111101001","111111111111110111","111111111111011101","111111111111110101","000000000000001001","000000000000000111","000000000000001010","111111111111101111","111111111111100000","111111111111100101","000000000000010000","000000000000010111","111111111111101000","000000000000011011","111111111111111100","111111111111101010","111111111111111101","000000000000000111","000000000000011011","111111111111010101","111111111111011110","111111111110111001","111111111111110010","111111111111101010","111111111111111101","111111111111111001","000000000000000111","111111111111111111","000000000000000111","111111111111100000","111111111111001011","111111111111011011","111111111111001100","111111111111111000","000000000000000000","111111111111011101","111111111111001001","111111111111110011","111111111111100110","111111111111110111","111111111111111011"),
("000000000000000110","000000000000110010","000000000000010100","111111111111110000","111111111111111100","111111111111111101","000000000000100000","111111111111011110","000000000000000100","111111111111111110","111111111111010000","111111111111010000","111111111111110100","000000000000001000","000000000000010000","111111111111110000","000000000000000110","111111111111111001","111111111111010000","111111111111111100","000000000000001001","000000000000100010","000000000000010011","000000000000001011","111111111111101101","000000000000010100","111111111111011101","000000000000001010","000000000000100010","111111111111101001","000000000000001000","111111111111100101","111111111111110011","111111111111101001","111111111111001110","000000000000001001","000000000000000110","111111111111110111","111111111111010000","111111111111101100","111111111111001010","111111111111010000","111111111111001011","111111111110110101","111111111111111010","000000000000010110","111111111111111001","000000000000101100","111111111111111111","111111111111110110","000000000000011100","000000000000000100","111111111111111001","111111111111100011","111111111111010101","000000000000011011","111111111111100111","000000000000010000","000000000000000000","111111111111101110","000000000000010110","000000000000001101","000000000000001010","000000000000001001","111111111111000011","000000000000010110","000000000000000011","000000000000000110","000000000000011011","111111111111101111","111111111111101011","111111111111010010","000000000000001101","000000000000010100","000000000000000100","111111111111011001","000000000000000001","111111111111101010","000000000000001010","000000000000100110","000000000000001011","000000000000000010","000000000000100010","000000000000001110","111111111111101101","111111111111110110","111111111110101010","111111111111100111","111111111111110011","111111111111110000","000000000000001001","111111111111101111","111111111111100100","000000000000001001","111111111111110100","111111111111001111","111111111111101001","000000000000100001","000000000000001010","000000000000001100","000000000000001000","111111111111011110","111111111111110111","111111111111101101","111111111111111000","111111111111111101","000000000000001000","111111111111100100","111111111110110110","111111111111110111","111111111111110011","111111111111110101","000000000000011010","111111111111111110","000000000000000000","000000000000000000","000000000000000100","111111111111000111","111111111111100000","111111111111010011","111111111111101111","111111111111101111","111111111111011010","111111111111100011","111111111111110000","000000000000000001","111111111111111111","111111111111100100"),
("000000000000100101","000000000000111101","000000000000010111","000000000000011010","000000000000000110","000000000000000001","000000000000110010","111111111111100100","000000000000000011","000000000000010000","111111111111010001","111111111111110101","000000000000000010","000000000000010100","000000000000010100","000000000000001011","000000000000100010","111111111111111101","111111111111011100","000000000000001011","000000000000001101","000000000000000101","000000000000001001","111111111111111110","111111111111110101","000000000000001110","111111111111010000","111111111111111111","111111111111111001","111111111111100100","000000000000001110","111111111111100111","111111111111011111","111111111111111111","111111111111011111","111111111111101110","000000000000001011","111111111111110110","111111111111011100","111111111111110111","111111111110110111","111111111111101110","111111111111011110","111111111111101010","000000000000000001","111111111111111001","111111111111110010","000000000000010111","111111111111110000","000000000000011001","000000000000100100","111111111111111010","000000000000010011","111111111111110000","111111111111010000","000000000000100000","111111111111110010","111111111111111011","000000000000000100","000000000000001100","111111111111100110","111111111111111000","000000000000010110","000000000000100000","111111111111100110","111111111111111011","111111111111111111","000000000000001101","000000000000111010","111111111111110000","000000000000000001","111111111111110101","111111111111110111","111111111111110001","000000000000000000","111111111111010101","000000000000000110","000000000000000000","000000000000001100","000000000000011001","000000000000000011","000000000000000111","000000000000010111","000000000000000000","111111111111110111","000000000000010101","111111111110111011","111111111111011111","000000000000001111","111111111111111001","000000000000001101","000000000000000110","111111111111111011","000000000000010011","111111111111111011","111111111111010100","111111111111101011","000000000000010101","111111111111110011","111111111111110001","000000000000101011","111111111111100000","111111111111110011","000000000000001011","111111111111111101","000000000000011110","111111111111111110","111111111111100100","111111111111010000","000000000000001011","000000000000001101","111111111111100110","000000000000010110","111111111111111011","111111111111111010","000000000000000000","000000000000011011","111111111111000000","111111111111010001","111111111110111111","000000000000010010","000000000000000010","111111111111001101","111111111110110101","000000000000000100","111111111111100010","000000000000011000","111111111111101110"),
("000000000000100011","000000000000100100","000000000000011000","000000000000000000","111111111111111100","000000000000001111","000000000000001111","111111111111100010","000000000000001011","111111111111101000","000000000000000010","000000000000000111","111111111111110010","000000000000111010","111111111111011011","000000000000000001","000000000000010101","111111111111111000","111111111111100101","111111111111100110","111111111111110110","111111111111101000","000000000000010010","000000000000000111","111111111111111100","111111111111111110","111111111111110000","111111111111111100","111111111111101011","111111111111110001","111111111111110110","111111111111101010","111111111111010101","111111111111010101","000000000000001010","111111111111100000","000000000000000101","111111111111111101","111111111111100010","111111111111101001","111111111110111011","000000000000001000","111111111111100110","000000000000011111","000000000000010110","000000000000000001","111111111111101101","111111111111111101","111111111111101000","111111111111110110","000000000001000011","000000000000010001","000000000000001011","111111111111010100","111111111111011011","111111111111111000","111111111111100110","111111111111111000","000000000000011001","000000000000001100","111111111111101110","000000000000001110","000000000000010110","000000000000011000","111111111111100100","000000000000001110","000000000000000101","000000000000001110","000000000000111111","111111111111101010","000000000000000000","111111111111110100","111111111111100110","111111111111101010","111111111111100110","111111111111000001","000000000000011110","111111111111101100","000000000000100001","000000000000010111","111111111111111001","000000000000000101","000000000000011110","000000000000000000","111111111111100100","000000000000001011","111111111110101100","111111111111110001","000000000000011110","111111111111110111","000000000000010110","111111111111101111","111111111111110111","000000000000001000","111111111111101100","111111111111011010","111111111111110110","000000000000000101","111111111111101000","111111111111111100","000000000000010110","111111111111101110","111111111111101000","111111111111110011","000000000000101000","000000000000101111","111111111111111100","111111111111100010","111111111111011000","000000000000001110","000000000000010000","111111111111110000","000000000000000101","111111111111100010","000000000000001101","000000000000000101","111111111111110001","111111111111100100","111111111111101010","111111111110111010","111111111111111101","000000000000011100","111111111111101101","111111111110011011","000000000000011100","111111111111111100","000000000000011110","111111111111101101"),
("000000000000010001","000000000000100000","000000000000010010","000000000000001111","111111111111111000","000000000000001100","000000000000011110","000000000000001110","000000000000001001","111111111111111011","000000000000001001","000000000000000000","111111111111111000","000000000000100100","111111111111100111","000000000000011110","000000000000010011","000000000000001101","000000000000000011","111111111111101101","000000000000001111","111111111111111110","000000000000011000","000000000000000100","000000000000000000","000000000000010000","111111111111110110","000000000000000000","111111111111010010","111111111111111101","000000000000010111","111111111111101011","111111111111100011","111111111111101011","000000000000001001","111111111111001111","111111111111110101","111111111111101011","000000000000000000","111111111111010111","111111111111011110","000000000000000010","000000000000011000","000000000000010111","111111111111111101","000000000000010101","000000000000100000","111111111111100101","111111111111101010","111111111111110010","000000000000100110","111111111111111110","000000000000001111","111111111111100001","111111111111000001","111111111111111011","111111111111110101","111111111111110011","111111111111111100","000000000000001011","111111111111111101","000000000000001010","000000000000001010","000000000000010110","111111111111110001","000000000000010100","111111111111111111","000000000000001011","000000000000100001","111111111111011100","000000000000011010","111111111111101010","111111111111101111","000000000000000010","111111111111010110","111111111110110011","000000000000000110","111111111111111100","111111111111100110","000000000000001101","000000000000011001","111111111111101110","000000000000011001","000000000000010100","111111111111100111","000000000000010010","111111111111010000","111111111111101111","000000000000001110","111111111111110101","000000000000000101","111111111111111111","111111111111111001","000000000000011110","111111111111110100","111111111111110101","111111111111011101","000000000000001010","111111111111100011","111111111111110111","000000000000011010","000000000000000000","000000000000000111","111111111111110010","000000000000100110","000000000000100111","111111111111111001","111111111111011001","111111111111100010","000000000000001010","000000000000000000","111111111111101111","000000000000010010","111111111111010101","000000000000000000","000000000000011100","000000000000000010","111111111111001101","111111111111101110","111111111111010001","000000000000000010","000000000000111011","000000000000001000","111111111101100000","000000000000001101","000000000000000000","000000000000011011","111111111111101011"),
("000000000000100110","000000000000000100","000000000000011010","000000000000000111","111111111111101101","000000000000010101","000000000000001011","111111111111111010","000000000000010001","111111111111101001","000000000000100010","000000000000001011","000000000000000001","000000000000011110","111111111111100010","111111111111111111","000000000000011010","111111111111111100","000000000000011100","000000000000000100","000000000000000010","000000000000001100","000000000000001101","000000000000011010","111111111111101111","000000000000010011","000000000000000100","000000000000010001","000000000000000100","000000000000000100","000000000000011000","000000000000001011","111111111111111010","000000000000001001","000000000000011100","111111111111011100","000000000000000011","000000000000000001","111111111111111110","111111111111101100","111111111111100110","111111111111111101","000000000000101001","111111111111111111","000000000000100101","111111111111111010","000000000001001100","111111111111100011","111111111111110011","111111111111110100","000000000000001010","000000000000011000","111111111111111001","111111111111101011","111111111111000111","000000000000001011","111111111111100110","111111111111101111","111111111111100111","000000000000000000","111111111111100110","000000000000000001","000000000000001011","000000000000010111","111111111111111001","000000000000000100","111111111111100101","000000000000001000","000000000000100100","111111111111101000","111111111111111001","111111111111110001","000000000000001001","111111111111100110","111111111110111110","111111111111000001","000000000000100010","111111111111110111","111111111111110001","000000000000000000","000000000000010011","000000000000000000","000000000000000000","000000000000011110","111111111111111011","111111111111111010","111111111110111101","111111111111101011","000000000000100010","111111111111110001","111111111111100110","000000000000000010","000000000000000101","000000000000000000","000000000000000010","000000000000000111","111111111110111111","111111111111111001","000000000000001001","111111111111100111","000000000000100010","111111111111111001","000000000000000111","111111111111110010","000000000000011101","000000000000011001","000000000000000100","000000000000011110","111111111111011101","111111111111111001","000000000000001101","111111111111111111","000000000000100011","111111111111011110","000000000000100110","000000000000010110","000000000000000011","111111111111100100","111111111111110001","111111111111001110","111111111111110101","000000000000110101","000000000000001000","111111111101100110","000000000000001011","000000000000011000","000000000000011000","111111111111011110"),
("000000000000000101","000000000000000110","000000000000001001","000000000000000000","111111111111111010","000000000000010100","111111111111111011","111111111111111100","000000000000001010","111111111111100110","000000000001000000","000000000000100001","000000000000001011","000000000000110000","111111111110110100","111111111111111010","000000000000000000","000000000000001001","000000000000011010","111111111111110010","000000000000000000","000000000000010001","111111111111111011","000000000000010000","111111111111111001","000000000000100011","000000000000001101","111111111111111110","111111111111111100","111111111111011010","111111111111110111","111111111111111001","000000000000010000","111111111111110010","000000000000010010","111111111111011111","111111111111101010","000000000000000110","000000000000001000","111111111111100010","111111111111000100","000000000000100111","000000000000111111","000000000000011110","000000000000001011","111111111111111011","000000000000101110","111111111111100100","000000000000000110","111111111111110000","111111111111011101","000000000000000100","111111111111100011","111111111111101010","111111111111101000","000000000000011011","000000000000000011","111111111111111011","111111111111101010","111111111111111101","111111111111101001","111111111111111101","111111111111110111","000000000000001110","111111111111111111","111111111111110101","111111111111011110","000000000000001000","000000000001000011","111111111111110011","000000000000010101","000000000000001000","111111111111111100","000000000000000111","111111111110111111","111111111110111011","000000000000001011","111111111111101110","111111111111101110","000000000000011111","000000000000000000","000000000000001001","000000000000011001","000000000000011101","111111111111110011","111111111111101101","111111111110101101","111111111111100010","000000000000100010","111111111111110111","111111111111100001","000000000000000110","111111111111110110","111111111111111101","000000000000001111","111111111111111100","111111111111000010","000000000000000001","111111111111101100","111111111111110111","000000000000100101","000000000000010100","111111111111111110","000000000000000101","000000000000100011","000000000000100111","000000000000000111","000000000000100110","000000000000000010","111111111111110100","000000000000000100","000000000000000000","000000000000000000","111111111111111011","000000000000101000","111111111111110011","111111111111111111","111111111111100111","111111111111111000","111111111111110001","000000000000001000","000000000000011011","000000000000001100","111111111110101000","000000000000010110","111111111111111010","000000000000011010","111111111111100111"),
("111111111111111001","111111111111100010","111111111111110101","000000000000011110","111111111111100101","000000000000010111","111111111111111010","111111111111110000","000000000000010101","111111111111100001","000000000000111011","000000000000010100","000000000000010000","000000000000111000","111111111111010100","111111111111110101","000000000000000011","000000000000001001","000000000000011011","111111111111111000","111111111111110111","111111111111111110","000000000000000000","000000000000001110","111111111111110000","000000000000100100","111111111111111101","000000000000001011","000000000000001011","111111111111110101","000000000000001001","000000000000000101","000000000000001110","111111111111111100","000000000000101010","111111111111101110","111111111111111000","000000000000100010","000000000000010001","111111111111110010","111111111110101011","000000000000100001","000000000000101001","111111111111110101","000000000000000010","000000000000000110","000000000000110101","000000000000010110","000000000000000101","000000000000010001","111111111110111111","000000000000000101","111111111111101100","111111111111111101","111111111111110110","000000000000001101","111111111111101100","111111111111101000","000000000000000000","111111111111110100","111111111111100100","000000000000000110","111111111111101101","000000000000000100","000000000000011111","111111111111101001","111111111111111011","111111111111101001","000000000000101101","111111111111111011","000000000000010000","000000000000000100","000000000000000011","111111111111111111","000000000000000000","111111111111010011","000000000000010001","111111111111111001","000000000000001101","000000000000001111","111111111111110001","000000000000000111","000000000000011110","000000000000101010","000000000000001001","111111111111100101","111111111110100100","111111111111011110","000000000000011001","000000000000100000","111111111111110010","111111111111011110","000000000000010110","000000000000001010","111111111111111010","000000000000001010","111111111111011001","000000000000001010","000000000000010000","000000000000010101","000000000000000111","000000000000110101","111111111111101101","000000000000001010","000000000000001010","000000000000001111","000000000000000000","000000000000011100","000000000000001110","111111111111111011","111111111111111111","111111111111100000","000000000000000100","111111111111111010","000000000000101110","111111111111101110","000000000000000000","111111111111100111","000000000000100100","111111111111101011","111111111111111111","111111111111110001","000000000000101101","111111111111111011","000000000000100010","000000000000000000","111111111111101010","111111111111110001"),
("000000000000010100","111111111111101001","000000000000001010","000000000000001011","111111111111110111","000000000000001101","000000000000001101","111111111111100110","000000000000010100","111111111111101111","000000000000011011","000000000000010001","000000000000100001","000000000000001000","000000000000011011","111111111111111000","111111111111111000","111111111111101101","000000000000100010","111111111111101101","111111111111110010","111111111111101111","111111111111110100","000000000000011010","111111111111110110","000000000000100000","111111111111111010","111111111111100111","000000000000010000","000000000000000001","000000000000010101","000000000000001101","111111111111011111","111111111111110110","000000000000001001","111111111111110100","000000000000000000","000000000000001010","000000000000001001","000000000000000010","111111111111010101","000000000000001000","111111111111110111","000000000000011001","000000000000000010","000000000000110010","000000000000001110","000000000000101011","000000000000000010","000000000000001010","111111111111001101","000000000000001011","111111111111111111","000000000000000001","111111111111110011","000000000000011100","111111111111111110","111111111111110110","000000000000000010","111111111111110000","111111111111100001","111111111111101100","111111111111111110","111111111111110001","000000000000001100","111111111111110111","000000000000010111","111111111111111111","000000000000001011","111111111111110101","111111111111110111","000000000000011000","000000000000000011","000000000000000111","111111111111101111","111111111111011000","000000000000000101","000000000000000010","000000000000100010","000000000000001100","000000000000001001","111111111111011101","000000000000101011","000000000000001100","111111111111101001","000000000000001001","111111111110111111","111111111111111001","000000000000010100","000000000000000111","000000000000110111","111111111111101000","111111111111110001","000000000000000000","111111111111111001","111111111111101010","111111111110111010","111111111111101001","000000000000001101","000000000000001000","111111111111101110","000000000000010011","111111111111110101","111111111111110001","111111111111111010","000000000000001100","000000000000000000","000000000000010111","000000000000000000","000000000000010110","000000000000001001","111111111111101000","111111111111110101","111111111111111010","000000000000001011","000000000000000101","000000000000001011","111111111111110000","000000000000000000","111111111111100100","111111111111100100","111111111111101101","000000000000001110","000000000000011111","000000000000011001","111111111111110010","111111111111110110","111111111111110011"),
("000000000000010101","111111111111011110","000000000000100011","111111111111111001","111111111111111100","000000000000001011","111111111111111111","111111111111100110","111111111111110111","111111111111101000","111111111111111100","111111111111110010","111111111111101011","000000000000010010","000000000000101000","111111111111100011","000000000000000010","000000000000001010","000000000000001101","000000000000000110","000000000000000101","111111111111010100","111111111111110111","111111111111111011","111111111111101011","000000000000001110","111111111111101111","111111111111110111","000000000000000001","000000000000000011","000000000000001010","111111111111110010","111111111111110001","000000000000000000","000000000000010000","111111111111110000","000000000000010011","000000000000001000","000000000000000011","111111111111111010","111111111111111110","000000000000001111","000000000000001001","111111111111111110","111111111111110100","000000000000011101","000000000000000000","000000000000010100","000000000000000000","000000000000001000","111111111111101101","000000000000000111","111111111111110000","111111111111110111","000000000000011001","000000000000100000","000000000000001101","111111111111110010","000000000000001111","111111111111101011","111111111111111101","111111111111111111","111111111111111101","111111111111111010","111111111111101111","000000000000001101","000000000000101010","111111111111111111","000000000000010111","111111111111110000","111111111111111111","111111111111110011","000000000000010010","000000000000001000","111111111111101111","111111111111110001","000000000000001111","000000000000001100","111111111111111100","000000000000001001","000000000000011010","111111111111111010","000000000000100111","000000000000000111","111111111111101110","000000000000110101","111111111111110010","111111111111101010","111111111111110111","000000000000000000","000000000000111100","111111111111100010","111111111111110100","111111111111110110","111111111111110111","000000000000100100","111111111111101101","111111111111110110","111111111111101000","111111111111111000","000000000000011101","000000000000100000","000000000000000011","111111111111110011","111111111111110001","000000000000001110","000000000000001101","000000000000100111","000000000000010110","000000000000111001","000000000000001001","111111111111001000","111111111111110011","111111111111110010","000000000000001010","111111111111110010","111111111111100000","111111111111101010","000000000000011011","111111111111111110","111111111111101101","111111111111111000","000000000000011100","000000000000101101","000000000000101010","111111111111101101","111111111111110010","111111111111110111"),
("111111111111100001","111111111111000100","000000000000011010","000000000000001110","000000000000011111","000000000000000000","000000000000011100","000000000000001101","111111111111111000","111111111111011110","000000000000000000","111111111111010100","111111111111110110","111111111111110110","000000000000111010","111111111111111110","000000000000001011","000000000000001110","000000000000010000","111111111111111111","111111111111100101","111111111111010110","000000000000000100","111111111111100000","000000000000000000","000000000000000101","000000000000000001","000000000000001111","111111111111101110","000000000000001111","111111111111100110","000000000000001000","000000000000000011","000000000000000110","000000000000000101","111111111111111011","000000000000011100","111111111111110101","000000000000001000","000000000000000100","111111111111110001","111111111111011011","000000000000000100","000000000000000101","000000000000010000","000000000000010001","000000000000011110","000000000000011010","111111111111111100","000000000000011000","111111111111100110","000000000000010010","111111111111111001","111111111111110010","000000000000001101","000000000000001111","000000000000100111","000000000000000000","000000000000011011","111111111111111111","111111111111110101","111111111111110011","111111111111101111","000000000000000110","111111111111101101","000000000000001011","000000000000010101","000000000000000000","000000000000010000","000000000000010100","111111111111110100","111111111111111000","000000000000001000","000000000000000000","111111111111111000","000000000000000001","000000000000010011","111111111111111011","000000000000010000","000000000000000001","111111111111111001","111111111111110001","000000000001001000","000000000000000011","111111111111110001","000000000000100111","000000000000010011","111111111111111001","111111111111111100","000000000000010000","000000000000100000","111111111111101011","000000000000010010","111111111111111010","000000000000011101","000000000000011010","000000000000011001","111111111111110000","000000000000001001","111111111111001100","111111111111111011","000000000000010100","111111111111111101","111111111111110000","111111111111101100","000000000000001011","111111111111111001","000000000000100101","000000000000000100","000000000000101100","111111111111111101","111111111111011000","000000000000001110","000000000000010011","000000000000100000","000000000000001010","000000000000000101","000000000000000101","000000000000000101","111111111111101111","111111111111011110","111111111111110011","111111111111110110","000000000000101100","000000000000010110","111111111111100111","111111111111110100","000000000000010100"),
("111111111111101011","111111111111100010","000000000000000111","111111111111101010","000000000000000000","000000000000000100","000000000000000111","000000000000000000","111111111111100110","111111111111110011","111111111111010011","111111111111101000","111111111111110101","111111111111110011","000000000000110001","111111111111100111","000000000000000100","111111111111110010","000000000000010110","000000000000010100","111111111111111011","000000000000001101","000000000000110000","111111111111011111","000000000000010110","111111111111111001","111111111111100101","111111111111110101","000000000000000111","000000000000010110","111111111111111100","111111111111111001","000000000000100001","111111111111111110","111111111111101010","111111111111110000","000000000000100100","000000000000010010","000000000000100010","000000000000000101","111111111111100110","111111111111101011","000000000000000100","111111111111101110","000000000000011100","111111111111110101","000000000000001101","000000000000010110","000000000000010011","000000000000010111","111111111111101011","000000000000001110","111111111111111111","000000000000011101","000000000000010010","000000000000000111","000000000000110000","000000000000011110","000000000000011111","000000000000000111","000000000000100001","111111111111100100","000000000000001100","111111111111111100","111111111111000101","000000000000011111","000000000000010110","111111111111111100","000000000000010001","111111111111111000","000000000000001101","111111111111111010","000000000000101010","000000000000010001","111111111111111110","000000000000000010","000000000000011000","000000000000001101","000000000000010000","000000000000010000","111111111111111000","000000000000100001","000000000000101000","111111111111111111","111111111111111010","000000000000101100","000000000000001111","111111111111111111","000000000000000001","000000000000001000","000000000000010001","111111111111111101","000000000000000110","000000000000000011","000000000000001011","000000000000000110","000000000000000000","000000000000010101","000000000000001001","111111111111011001","000000000000001001","111111111111110001","111111111111111110","000000000000000001","111111111111111110","000000000000000111","111111111111110011","000000000000000111","000000000000000101","000000000000011100","111111111111110001","111111111111100110","000000000000000010","000000000000000010","000000000000011101","111111111111111111","000000000000000001","000000000000000100","000000000000000000","000000000000001111","111111111111110000","000000000000001100","111111111111101111","000000000000001111","000000000000100010","111111111111110010","111111111111101100","000000000000010001"),
("111111111111011001","000000000000001001","111111111111111111","111111111111011111","111111111111111011","111111111111110100","111111111111111011","000000000000010111","111111111111111001","000000000000000101","111111111111111100","111111111111100110","000000000000000111","111111111111010110","000000000000111001","111111111111111101","000000000000000111","111111111111110010","111111111111111100","111111111111111000","111111111111111111","000000000000000010","000000000000010110","111111111111101010","000000000000001001","000000000000001011","111111111111110000","111111111111110111","111111111111110100","000000000000100111","000000000000000100","000000000000000000","111111111111111100","111111111111111100","111111111111100111","111111111111110111","111111111111111110","111111111111111110","111111111111111110","000000000000100010","111111111111111111","111111111111110000","000000000000001010","111111111111101110","000000000000000111","111111111111110111","111111111111110101","000000000000100101","000000000000011100","000000000000000101","111111111111101111","000000000000000001","000000000000001010","000000000000001110","111111111111111110","000000000000011111","000000000000011001","000000000000010010","111111111111111111","000000000000000110","000000000000001110","111111111111101001","111111111111101011","111111111111111001","111111111110111101","111111111111111111","111111111111111110","000000000000001011","000000000000010110","000000000000011010","111111111111101110","111111111111101001","000000000000000010","111111111111110010","000000000000001101","000000000000100101","000000000000000000","000000000000000000","000000000000010110","000000000000010000","111111111111101101","111111111111110110","000000000000111110","000000000000100101","111111111111101111","000000000000010111","000000000000100111","000000000000001010","111111111111111110","111111111111111101","000000000000100001","000000000000000110","111111111111110110","000000000000000000","111111111111101101","000000000000010111","000000000000000101","000000000000010001","000000000000100011","111111111111110010","000000000000000000","111111111111110010","000000000000010110","111111111111011110","111111111111111111","111111111111111101","000000000000000011","111111111111101110","111111111111110100","000000000000010111","111111111111111111","000000000000010111","000000000000010111","111111111111111000","000000000000000010","000000000000000010","000000000000000000","000000000000000110","111111111111101010","111111111111101110","111111111111111010","000000000000000000","111111111111110001","000000000000011001","000000000000110011","000000000000001000","111111111111110110","111111111111101111"),
("111111111111101111","000000000000100001","111111111111110101","111111111111001100","000000000000000000","111111111111110101","111111111111110011","000000000000101110","111111111111011110","000000000000010000","111111111111110011","000000000000000001","000000000000000101","111111111111101011","000000000000000101","000000000000000110","111111111111110101","111111111111010000","000000000000000110","000000000000010001","000000000000000000","000000000000001111","000000000000100111","111111111111101111","111111111111110011","000000000000001101","111111111111100000","111111111111011010","000000000000001100","111111111111101011","111111111111110000","111111111111111100","000000000000000000","111111111111101100","111111111111011111","111111111111111011","000000000000000000","111111111111110011","111111111111110111","000000000000000111","111111111111111011","000000000000001100","000000000000001101","000000000000000000","000000000000010101","111111111111111011","111111111111111011","000000000000001111","000000000000001000","000000000000000100","000000000000001001","111111111111110001","111111111111111000","000000000000001011","000000000000000001","000000000000000001","000000000000001100","111111111111111011","000000000000001110","111111111111101110","000000000000011101","111111111111111101","111111111111100010","111111111111111000","111111111110100100","111111111111101111","111111111111001001","111111111111111110","000000000000011100","111111111111110100","111111111111111110","111111111111111101","000000000000010010","111111111111110110","000000000000011010","000000000000001100","000000000000010111","111111111111110001","000000000000001111","000000000000001111","111111111111011110","000000000000000000","000000000000010101","000000000000101101","000000000000010100","111111111111110010","111111111111110010","000000000000011001","000000000000000100","111111111111110110","000000000000001010","000000000000000111","000000000000000000","000000000000001010","111111111111111001","111111111111010000","000000000000010101","111111111111111110","000000000000101110","000000000000000101","111111111111111111","000000000000001001","111111111111110111","000000000000001000","000000000000000000","000000000000001010","111111111111101111","111111111111110111","111111111111110101","111111111111110100","111111111111110100","000000000000010111","000000000000001011","000000000000001011","000000000000000100","111111111111110101","000000000000011010","000000000000001001","111111111111101110","000000000000001001","111111111111111011","000000000000001101","111111111111100110","000000000000010110","000000000000011101","111111111111111010","111111111111100000","111111111111110000"),
("000000000000000111","000000000000001011","111111111111111010","111111111111001011","000000000000001100","111111111111110000","111111111111110010","000000000000011011","111111111111101110","000000000000001010","111111111111100110","000000000000010001","111111111111111011","000000000000001010","000000000000000011","111111111111110001","111111111111110001","111111111111110101","000000000000001101","111111111111110010","111111111111111111","000000000000001111","000000000000010100","000000000000001110","000000000000000101","111111111111101100","111111111111010010","111111111111011001","111111111111111010","111111111111111110","000000000000000111","111111111111111001","000000000000010001","000000000000011000","111111111111110001","111111111111110100","000000000000000011","111111111111111011","111111111111011010","000000000000100111","111111111111101100","000000000000001010","000000000000001001","111111111111111100","000000000000010111","111111111111110100","000000000000001101","000000000000001011","000000000000100001","111111111111100000","000000000000000011","000000000000000000","000000000000100000","111111111111111001","000000000000000110","000000000000000001","000000000000000100","000000000000001000","000000000000001000","111111111111111010","111111111111101110","111111111111100010","111111111111011101","111111111111100011","111111111111001101","000000000000001000","111111111111011010","111111111111111100","111111111111111100","000000000000001001","111111111111111111","000000000000001110","111111111111110100","000000000000001101","000000000000000001","000000000000100100","000000000000001111","111111111111101010","111111111111110100","111111111111111011","111111111111110010","111111111111101110","000000000000101011","000000000000001001","111111111111101110","111111111111100001","111111111111110110","000000000000000000","111111111111111001","000000000000001100","000000000000000110","111111111111111101","111111111111101001","111111111111111011","111111111111110001","111111111111000011","111111111111111001","000000000000010000","000000000000100110","111111111111111100","000000000000010001","000000000000000011","111111111111100011","111111111111100011","111111111111101110","111111111111110100","111111111111110011","111111111111100101","111111111111010111","000000000000011110","111111111111100111","111111111111101110","000000000000001100","111111111111110110","111111111111101001","111111111111110110","111111111111111111","000000000000011011","111111111111001111","000000000000000110","000000000000011011","000000000000001001","111111111111111100","000000000000011010","000000000000000011","000000000000001100","111111111111110011","000000000000000011"),
("111111111111110010","000000000000100000","000000000000000011","111111111111100100","000000000000100111","000000000000001001","000000000000000011","000000000000001010","000000000000000111","000000000000011101","111111111111111111","000000000000010100","111111111111101100","000000000000001011","000000000000001001","111111111111111001","000000000000001100","000000000000001010","111111111111110010","111111111111111011","000000000000000101","111111111111111110","000000000000000101","111111111111101100","111111111111101100","000000000000000010","111111111111110010","111111111111100101","000000000000000000","111111111111100111","111111111111110111","111111111111111100","000000000000000011","111111111111111110","000000000000001001","111111111111111001","000000000000000110","000000000000010010","111111111111110111","000000000000001001","000000000000001010","000000000000110001","000000000000001101","111111111111110011","000000000000001111","111111111111110101","000000000000000111","111111111111111010","000000000000011011","111111111111100000","000000000000001100","000000000000010001","000000000000001110","000000000000010101","000000000000001111","000000000000000100","111111111111011111","111111111111100000","111111111111110011","111111111111101111","111111111111100101","111111111111011111","111111111111101011","000000000000000000","000000000000010011","000000000000000000","111111111110011111","111111111111111110","000000000000010000","000000000000000000","000000000000000101","111111111111101111","111111111111000110","000000000000001110","000000000000011011","000000000000110010","000000000000000010","111111111111011111","000000000000010100","000000000000100000","111111111111111110","111111111111101101","000000000000101111","111111111111011111","111111111111110110","111111111111100001","000000000000010100","000000000000110010","111111111111111001","000000000000001010","111111111111101010","111111111111100111","111111111111110010","000000000000001101","111111111111101010","111111111111001110","000000000000001000","000000000000000100","000000000000001011","111111111111110111","111111111111111111","000000000000000001","111111111111100011","111111111111111000","000000000000011111","111111111111110100","111111111111100101","111111111111110010","111111111111111110","000000000000010000","000000000000001010","111111111111101010","000000000000001000","000000000000011010","000000000000000010","111111111111100111","000000000000001010","000000000000001110","111111111111110010","000000000000001010","000000000000000001","000000000000010110","111111111111100111","000000000000011011","000000000000100010","000000000000001101","111111111111111001","111111111111110010"),
("111111111111111110","000000000000111111","111111111111110100","000000000000000010","000000000000000000","000000000000010010","111111111111111000","111111111111111001","111111111111111010","000000000000001101","111111111111111101","000000000000101111","111111111111101000","111111111111101110","111111111111111100","000000000000001100","000000000000001001","111111111111110110","111111111111101101","000000000000010011","111111111111111011","000000000000000000","000000000000000011","111111111111111111","000000000000000000","111111111111111011","111111111111110110","111111111111111011","111111111111110011","111111111111101010","111111111111110001","111111111111111111","000000000000001001","111111111111111101","111111111111101011","000000000000000110","111111111111111100","000000000000001001","111111111111011001","000000000000000000","000000000000010111","000000000000000011","000000000000001110","111111111111001101","111111111111110100","000000000000001110","000000000000001100","000000000000000011","000000000000011101","111111111111101010","000000000000001101","111111111111100111","000000000000010001","000000000000000001","000000000000000101","111111111111110110","111111111111010100","000000000000000001","000000000000001010","111111111111110011","111111111111010011","111111111111010100","000000000000000100","111111111111101110","000000000000000000","000000000000001100","111111111110110101","000000000000001101","000000000000110101","111111111111100101","111111111111101101","111111111111100110","111111111110110011","000000000000000110","000000000000010011","000000000000100010","000000000000001010","111111111111111101","111111111111101101","000000000000001100","111111111111011111","111111111111010111","000000000000001111","111111111111100010","000000000000000110","111111111111111100","111111111111110101","000000000000101101","000000000000001001","000000000000100100","000000000000001100","111111111111111111","000000000000001000","000000000000010101","111111111111100011","111111111111100001","111111111111100101","111111111111111000","111111111111011101","111111111111011101","000000000000010011","111111111111111010","111111111111011111","111111111111101001","000000000000010110","000000000000000100","111111111111111110","111111111111110000","111111111111100101","111111111111111111","000000000000001011","111111111111011101","000000000000011010","000000000000001000","111111111111111111","111111111111110101","000000000000000000","000000000000000011","111111111111010100","111111111111111011","000000000000000000","000000000000001000","111111111111110110","000000000000010110","000000000000100010","111111111111111000","111111111111111010","111111111111100010"),
("111111111111101001","000000000000010100","000000000000001111","111111111111110101","000000000000001101","000000000000001100","111111111111101001","111111111111101110","000000000000010100","000000000000011101","111111111111111111","000000000000111110","111111111111101010","000000000000000110","111111111111110101","000000000000001111","000000000000001010","000000000000000100","111111111111101110","111111111111110011","000000000000001101","111111111111110100","000000000000000010","111111111111111000","111111111111110101","111111111111101111","000000000000010000","111111111111101101","111111111111110011","111111111111111010","111111111111110010","111111111111011101","111111111111100001","111111111111001100","111111111111110100","111111111111111011","000000000000001010","111111111111110001","111111111111100000","000000000000010001","111111111111111011","111111111111111100","111111111111111100","111111111111011000","000000000000001001","000000000000001010","000000000000001001","000000000000100110","000000000000000000","111111111111111111","000000000000100000","111111111111101010","000000000000010011","111111111111110011","000000000000011000","111111111111110100","111111111111011110","000000000000000101","111111111111101110","111111111111111110","111111111111101001","111111111111010101","000000000000001011","111111111111110010","000000000000001010","000000000000000010","111111111111110111","111111111111111101","000000000000101101","111111111111100111","000000000000000000","111111111111100011","111111111111000011","000000000000001101","111111111111111000","000000000000010111","111111111111110101","111111111111101100","111111111111111000","000000000000010001","111111111111101001","111111111111010011","000000000000010000","111111111111011010","000000000000001000","111111111111101011","111111111111110100","000000000000011100","000000000000000100","000000000000010011","111111111111111110","000000000000101001","111111111111111100","000000000000000000","111111111111101100","111111111111101001","000000000000011101","111111111111110110","111111111111010110","111111111111111101","111111111111100101","000000000000001010","111111111111111000","000000000000001000","000000000000000011","000000000000000101","111111111111111000","000000000000001010","111111111111110000","111111111111100010","000000000000001100","111111111111010101","000000000000011101","000000000000011010","000000000000000010","111111111111110011","111111111111111001","111111111111110000","111111111111101100","000000000000001000","111111111111101010","111111111111101110","000000000000010001","111111111111110001","111111111111111100","111111111111100101","000000000000000101","111111111111101000"),
("111111111111011001","000000000000100000","111111111111100100","000000000000001001","000000000000001010","111111111111110011","000000000000011000","111111111111110001","000000000000001000","000000000000001100","000000000000001010","000000000000100101","111111111111101101","111111111111111110","111111111111101100","000000000000000001","111111111111111000","000000000000010010","111111111111111111","000000000000001000","000000000000110111","000000000000001000","111111111111110001","111111111111111001","000000000000000000","111111111111101001","111111111111110101","111111111111101101","000000000000101001","111111111111101110","111111111111111100","111111111111101001","111111111111100110","111111111111101110","111111111111111110","000000000000001010","111111111111111110","000000000000000000","111111111111011111","000000000000010001","111111111111110111","000000000000010000","000000000000010011","111111111111111000","111111111111100011","111111111111101110","000000000000010001","000000000000100000","111111111111101111","111111111111111001","000000000000010101","111111111111111111","000000000000000011","111111111111110000","000000000000101111","111111111111111100","111111111111110010","111111111111111110","000000000000010011","000000000000010011","111111111111010101","111111111111100100","000000000000001110","111111111111111110","111111111111111000","000000000000001110","111111111111110110","111111111111100001","000000000000010010","111111111111100110","111111111111110110","111111111111101001","111111111111100010","000000000000010111","000000000000001000","000000000000010100","111111111111101000","111111111111011100","000000000000001100","000000000000011000","111111111111111000","111111111111010111","000000000000000000","111111111111101010","111111111111111010","111111111111001001","111111111111111010","000000000000010100","111111111111110011","000000000000000011","000000000000001001","111111111111110111","000000000000010111","000000000000000101","000000000000001111","111111111111100101","000000000000000011","111111111111101000","111111111111011001","111111111111010000","111111111111111110","000000000000000100","111111111111001110","000000000000010011","000000000000100110","000000000000001100","111111111111100100","000000000000000100","111111111111110011","111111111111101111","111111111111101100","111111111111110000","111111111111111111","111111111111111110","111111111111010111","111111111111110111","111111111111111011","000000000000011000","111111111111010110","111111111111100101","000000000000000000","000000000000000011","000000000000011101","000000000000011011","000000000000010011","000000000000000111","111111111111110000","111111111111010101"),
("000000000000001100","111111111111101010","111111111111100110","000000000000010010","111111111111101111","000000000000101001","000000000000100101","111111111111110011","000000000000001111","000000000000000011","000000000000110011","111111111111101011","000000000000010000","111111111111110001","111111111111111001","000000000000100110","000000000000011001","111111111111111011","000000000000000000","111111111111111111","000000000000011011","111111111111110001","000000000000001111","111111111111111001","111111111111100010","000000000000011011","111111111111011110","000000000000001110","000000000000011110","111111111111010100","000000000000011100","111111111111101011","000000000000010010","111111111111011010","000000000000011101","111111111111000110","000000000000101111","111111111111101001","111111111111110001","111111111111110010","111111111111011000","111111111111111111","000000000001011101","000000000000111011","111111111111011001","111111111111000111","000000000000011100","000000000000110101","111111111110111011","111111111111101000","111111111111101010","111111111111101001","111111111111100111","111111111111110111","000000000000111110","000000000000000111","111111111111111000","000000000000011101","111111111111100111","000000000000010001","111111111111001000","000000000000010110","000000000000100001","111111111111111101","000000000000001110","111111111111110001","000000000000011100","111111111111110011","000000000000000011","111111111111111000","111111111111110010","111111111111101111","000000000000001010","000000000000100100","111111111111101000","111111111111111111","000000000000101001","000000000000000011","000000000000101011","000000000000001000","111111111111110101","111111111111101010","000000000000100001","000000000000000101","111111111111101011","111111111111001000","000000000000100111","111111111111110000","111111111111111011","111111111111101000","111111111111100010","111111111110110100","000000000000000001","000000000000011010","111111111111100011","000000000000000010","111111111111111000","000000000000101000","111111111111000110","000000000000000111","000000000000011101","000000000000001011","111111111111011000","111111111111100100","000000000000010110","000000000000100101","111111111111010000","000000000000001010","111111111111110010","111111111111110111","111111111111001001","000000000000010111","111111111111111101","111111111110111111","111111111111001010","000000000000000101","000000000000001101","000000000000111110","111111111111110111","111111111111101110","000000000001000111","000000000000110111","000000000000111101","000000000000000101","000000000000110110","111111111111110110","000000000000010001","111111111111010100"),
("000000000000100011","111111111111001000","111111111111011010","111111111111111001","000000000000101011","111111111111111000","000000000000001001","000000000000011100","000000000000010101","111111111111100111","000000000000101010","111111111111100001","000000000000100010","000000000000001110","111111111111101100","000000000000000110","000000000000010000","000000000000001110","111111111111101100","000000000000001100","000000000000011001","000000000000001000","000000000000001111","111111111111111010","111111111111011101","111111111111110100","111111111111110011","000000000000011010","000000000000010100","000000000000000101","000000000000010101","111111111111100100","111111111111110111","111111111111100011","000000000000111111","000000000000000000","000000000000010001","000000000000000100","000000000000000010","000000000000010100","111111111111110011","000000000000000010","000000000000001110","000000000000011100","111111111111100000","000000000000000001","000000000000000010","111111111111111011","111111111111101010","111111111111101101","111111111111110110","000000000000001001","111111111111011110","000000000000001100","000000000000011011","000000000000100110","000000000000001001","000000000000011110","000000000000000100","111111111111110000","111111111111110011","000000000000010001","000000000000000110","111111111111111101","000000000000011100","111111111111110000","000000000000001110","111111111111100001","000000000000001000","111111111111101111","111111111111110010","000000000000000000","000000000000010111","000000000000010001","111111111111110010","111111111111110100","000000000000001001","000000000000000011","000000000000000100","000000000000010101","111111111111100011","111111111111100011","000000000000001000","000000000000001010","111111111111110100","111111111111100010","000000000000000101","111111111111111001","111111111111011001","111111111111111010","111111111111001101","111111111111000000","111111111111010000","000000000000000100","111111111111110111","111111111111100110","000000000000000100","111111111111111011","000000000000000000","000000000000000100","000000000000001001","111111111111011111","111111111111010110","111111111111101010","000000000000001100","111111111111110011","000000000000001010","000000000000010001","111111111111101010","000000000000001001","111111111111110110","000000000000011011","111111111111011111","111111111111111111","111111111111101100","000000000000000111","111111111111001100","000000000000110010","000000000000010000","000000000000000110","000000000000001110","000000000000010101","000000000000000100","000000000000001000","000000000000000011","111111111111100110","000000000000011000","111111111111111110"),
("111111111111111111","111111111111000011","111111111111101110","000000000000001011","111111111111010101","000000000000000000","000000000000100100","000000000000001101","000000000000001000","000000000000001010","000000000000100110","111111111111110010","000000000000011101","111111111111111111","111111111111100110","000000000000011000","000000000000001111","000000000000111100","111111111111000100","000000000000011011","000000000000011010","111111111111110011","111111111111110011","000000000000000010","000000000000010110","000000000000010000","111111111111110001","000000000000000111","111111111111110000","111111111111110110","000000000000100000","111111111111010110","000000000000011101","111111111111101000","000000000000010110","111111111111111011","000000000000001010","000000000000101001","111111111111100110","111111111111011100","111111111111101110","111111111111110001","000000000000100101","000000000000101001","000000000000001001","111111111111011110","000000000000100000","111111111111100111","111111111111010011","111111111111011110","000000000000011111","000000000000110110","000000000000010111","000000000000000101","000000000000011010","111111111111100011","111111111111100000","000000000000000010","111111111111110111","111111111111110111","000000000000010110","000000000000001111","000000000000110111","111111111111100100","111111111111110010","000000000000000010","000000000000100011","000000000000000111","000000000000010001","111111111111100101","000000000000001010","000000000000101010","000000000000011000","000000000000100100","111111111111100101","111111111111100000","000000000000000100","000000000000001001","111111111111001110","111111111111110101","111111111111011001","000000000000011011","000000000000100001","111111111111101000","000000000000001101","111111111111110001","111111111111110000","111111111111100001","111111111111100010","111111111111011000","111111111111001011","111111111111110111","111111111111110010","000000000000011010","000000000000000000","111111111111101000","000000000000011000","111111111111111011","111111111111010111","111111111111111001","000000000000011000","111111111111100100","000000000000010011","000000000000010101","111111111111111111","000000000000100001","111111111111010010","111111111111101100","111111111111100111","000000000000010101","111111111111011010","000000000000011101","111111111111110010","111111111111100100","000000000000000111","000000000000010010","000000000000010010","000000000000011100","111111111111111011","000000000000010111","000000000000010101","000000000000101001","000000000000111101","000000000000001110","000000000000010000","111111111111111001","000000000000010001","111111111111100110"),
("111111111111111111","000000000000000111","111111111111110110","000000000000001100","111111111111110111","111111111111100101","000000000000000000","111111111111111011","000000000000010110","000000000000000001","000000000000001001","111111111111110011","000000000000001111","000000000000010101","000000000000101000","000000000000001011","111111111111011010","111111111111101100","111111111111101111","000000000000011110","000000000000100100","000000000000001110","111111111111110000","000000000000000010","000000000000011001","111111111111100111","111111111111110010","000000000000000101","000000000000001101","111111111111111011","111111111111111100","000000000000000100","111111111111101011","111111111111111001","000000000000011101","111111111111011101","000000000000011001","111111111111110010","111111111111100010","000000000000011100","111111111111111100","111111111111111111","000000000000000101","000000000000011011","111111111111111110","111111111111110111","111111111111101110","111111111111110011","000000000000001011","000000000000010101","000000000000001000","111111111111100110","000000000000010001","111111111111110101","000000000000011111","000000000000010000","000000000000000010","000000000000010010","000000000000001000","111111111111110101","000000000000001100","111111111111110100","000000000000100100","111111111111111101","111111111111111111","000000000000010101","111111111111110011","000000000000000010","000000000000001101","000000000000000001","000000000000000010","111111111111101101","000000000000101011","000000000000101001","000000000000100000","111111111111111011","111111111111100111","000000000000011001","000000000000010011","111111111111111011","111111111111111000","111111111111101000","000000000000000000","111111111111110010","111111111111111011","111111111111110011","000000000000000101","111111111111100110","111111111111111000","000000000000000101","111111111111100000","111111111111111100","000000000000011110","111111111111111111","000000000000100000","111111111111111111","111111111111110000","000000000000001110","111111111111100001","000000000000010111","111111111111110001","111111111111100100","111111111111100101","111111111111101101","111111111111111111","111111111111010101","000000000000001000","111111111111111101","111111111111011111","111111111111110000","000000000000000111","000000000000000000","111111111111101100","111111111111110101","111111111111111010","000000000000001100","000000000000010101","000000000000011101","111111111111111110","111111111111111110","111111111111101110","000000000000001101","000000000000001111","000000000000011101","000000000000000000","111111111111111000","000000000000000110","111111111111111010"),
("000000000000000101","111111111111110000","000000000000000010","000000000000001100","000000000000001010","111111111111110101","000000000000000100","000000000000010001","000000000000000000","111111111111111100","000000000000001110","000000000000001100","111111111111101110","000000000000001010","111111111111101010","111111111111101111","111111111111111100","111111111111111110","000000000000000001","000000000000000101","111111111111110101","000000000000001100","000000000000011101","111111111111110111","111111111111111000","000000000000010000","111111111111111100","000000000000001010","000000000000100000","000000000000000000","000000000000000000","000000000000011011","111111111111110011","000000000000000101","111111111111101100","000000000000010011","111111111111101100","000000000000000000","000000000000000100","111111111111111101","000000000000010000","000000000000000011","000000000000000001","000000000000000100","111111111111111011","000000000000011011","111111111111110101","111111111111100000","000000000000001000","111111111111111000","000000000000010000","000000000000000010","111111111111100111","000000000000001101","000000000000100001","111111111111110000","000000000000000110","000000000000001010","000000000000001000","000000000000000101","111111111111110110","000000000000011111","000000000000010001","111111111111110010","000000000000000110","111111111111101101","111111111111110110","111111111111111000","111111111111111111","111111111111111101","111111111111111111","111111111111111011","111111111111110110","000000000000100001","000000000000000011","000000000000011001","111111111111011110","000000000000011110","111111111111100011","111111111111111101","000000000000000010","000000000000001000","000000000000000101","000000000000000001","000000000000100010","111111111111101111","111111111111111010","000000000000000001","000000000000000010","000000000000000011","111111111111110001","111111111111111110","111111111111101010","111111111111111001","111111111111101100","000000000000010000","000000000000000001","000000000000000000","111111111111110110","000000000000011011","111111111111100010","111111111111110000","000000000000011110","000000000000001001","111111111111110101","111111111111101110","000000000000010000","000000000000000101","000000000000010100","111111111111110011","000000000000000000","111111111111111000","000000000000010110","000000000000010001","000000000000011101","000000000000011110","000000000000000110","111111111111111000","000000000000000010","000000000000000100","111111111111111011","111111111111100000","111111111111111100","111111111111101101","111111111111110101","111111111111110101","111111111111101010","000000000000001011"),
("000000000000000100","111111111111111011","000000000000100000","111111111111100101","000000000000011000","000000000000000000","111111111111100001","111111111111111111","000000000000100101","000000000000011101","111111111111011101","000000000000001101","111111111111111101","111111111111111101","000000000000011100","111111111111111011","000000000000011000","000000000000000101","000000000000001010","000000000000001001","111111111111011100","000000000000000011","000000000000100001","111111111111010101","111111111111101101","111111111111101110","111111111111111100","111111111111110000","000000000000111100","000000000000011101","111111111111011011","000000000000001111","111111111111110101","111111111111101000","111111111111111101","000000000000010001","000000000000000000","000000000000010101","000000000000000111","000000000000000000","000000000000000000","111111111111110111","111111111111111110","000000000000001110","000000000000001100","111111111111110110","000000000000011001","111111111111110001","000000000000000000","000000000000011100","000000000000010000","000000000000011100","111111111111100110","111111111111111000","000000000000001100","000000000000011010","000000000000001000","111111111111111011","111111111111101001","000000000000001000","111111111111110000","111111111111101111","111111111111101001","000000000000011000","111111111111101001","111111111111011011","111111111111101001","111111111111101010","000000000000000100","000000000000000010","111111111111111100","000000000000000111","111111111111100010","111111111111111110","000000000000010001","000000000000100100","111111111111100101","111111111111110111","000000000000010010","000000000000010101","111111111111110111","111111111111110111","111111111111111001","000000000000010011","000000000000010000","000000000000011011","000000000000010000","000000000000010010","000000000000000000","000000000000011110","000000000000001101","111111111111111000","000000000000010011","111111111111101101","111111111111101111","111111111111111110","000000000000000100","000000000000000010","000000000000000101","000000000000000011","000000000000000100","111111111111010001","111111111111101111","111111111111111011","000000000000000011","111111111111101101","000000000000010000","000000000000001000","000000000000011011","000000000000000111","111111111111111111","111111111111100000","000000000000010110","000000000000000000","000000000000010010","111111111111111001","111111111111110011","000000000000011100","111111111111100111","000000000000100101","111111111111100011","111111111111111110","111111111111111000","000000000000010010","000000000000010111","111111111111011011","111111111111010011","000000000000010111"),
("000000000000010100","111111111111111110","111111111111011110","000000000000010010","000000000000000101","000000000000010001","111111111111011000","000000000000001000","000000000000100100","111111111111101111","111111111111001010","111111111111111001","111111111111110100","111111111111010011","111111111111100101","111111111111101001","000000000000100000","111111111111111010","000000000000010011","000000000000100111","111111111111101011","111111111111001010","000000000000000100","111111111111010110","111111111111011010","000000000000110000","111111111111111010","000000000000010100","000000000000010011","000000000000000100","000000000000010111","000000000000100100","000000000000011011","111111111111111010","111111111111101001","111111111111110011","111111111111100100","000000000001001010","111111111111110001","000000000000100111","000000000000100111","000000000000011101","111111111111101100","111111111111011110","000000000000111011","000000000000010011","000000000000011011","111111111111111101","000000000000000001","000000000000000001","000000000000010000","000000000000100100","111111111111000000","000000000000011110","000000000000101000","000000000000001011","111111111111101101","000000000000000001","111111111111011000","000000000000000001","000000000000010000","000000000000101011","000000000000001111","111111111111100010","000000000000001001","111111111111100001","111111111111000110","111111111111111011","111111111111011110","111111111111011011","000000000000100110","000000000000100101","111111111111011001","111111111111101001","000000000000110101","000000000000010011","111111111111100111","000000000000010000","111111111111110011","000000000000011100","111111111111100101","000000000000011000","000000000000100110","111111111111101001","000000000000001100","111111111111100000","111111111111110110","000000000000110110","111111111111110110","111111111111111110","000000000000001100","111111111111110111","111111111111100101","111111111111110100","111111111110111111","111111111111110101","000000000000001110","000000000000111001","000000000000011001","111111111111111110","111111111111111111","111111111111111101","111111111111110110","111111111111110101","111111111111010101","111111111111111010","111111111111001011","111111111111100001","111111111111101100","111111111111100000","111111111111100111","000000000000000011","000000000000101010","000000000000100110","000000000000011100","000000000000010000","000000000000101000","000000000000011110","000000000000000000","000000000000101111","000000000000010110","111111111111010101","111111111111110011","111111111111011011","000000000000010000","111111111111010111","111111111111101011","000000000000000001"),
("000000000000000010","111111111111110100","111111111111010010","000000000000001001","000000000000000110","000000000000000100","111111111111101001","000000000000000011","111111111111111101","111111111111111011","111111111110111011","111111111111011100","111111111111101100","111111111111000100","111111111111111001","000000000000010001","000000000000001110","000000000000000111","000000000000000010","000000000000100000","111111111111100110","000000000000001001","111111111111110100","111111111111100100","111111111111111011","111111111111110100","111111111111111011","000000000000000000","000000000000001100","000000000000010000","000000000000001100","111111111111110100","000000000000010100","000000000000000110","111111111111110011","111111111111101110","111111111111111111","000000000000111000","111111111111010010","000000000000101001","000000000000010001","000000000000000111","000000000000000000","111111111111110100","000000000000001001","000000000000000001","000000000000001110","000000000000010000","111111111111110101","000000000000000000","111111111111110100","000000000000101101","111111111111110100","000000000000000000","000000000000001101","000000000000010001","111111111111101100","111111111111110011","111111111111111001","111111111111111111","000000000000000010","111111111111111010","000000000000011100","111111111111011101","111111111111110011","000000000000000001","000000000000000011","111111111111111101","111111111111010100","000000000000011110","111111111111101110","111111111111111101","111111111111110100","111111111111010100","000000000000010010","111111111111010000","000000000000001011","111111111111111011","111111111111111011","000000000000100000","111111111111101010","000000000000010111","000000000000011100","111111111111101011","000000000000000001","111111111111110111","000000000000001000","000000000000010110","111111111111110111","000000000000001101","000000000000000101","111111111111100100","111111111111110001","111111111111100010","111111111111011111","000000000000000010","000000000000010010","000000000000011001","000000000000100010","111111111111011001","000000000000010101","111111111111010110","111111111111111101","000000000000000100","000000000000000100","111111111111110101","111111111111100101","111111111111100110","111111111111010011","000000000000010010","111111111111101001","111111111111101110","111111111111110010","000000000000010001","000000000000011001","111111111111100101","111111111111110100","000000000000001111","111111111111101111","000000000000011101","000000000000010010","000000000000000010","111111111111111010","111111111111001110","000000000000100001","111111111111101101","000000000000001111","111111111111110001"),
("111111111111111101","111111111111111011","111111111111110110","111111111111111110","000000000000010001","000000000000000000","000000000000000000","000000000000000000","000000000000010011","000000000000000000","111111111110110010","111111111111011011","111111111111110000","111111111111100100","111111111111111000","000000000000000001","111111111111110011","000000000000001011","111111111111110000","111111111111111110","111111111111110111","000000000000001100","111111111111110000","111111111111011011","111111111111111000","000000000000000000","111111111111100100","000000000000100000","000000000000000111","111111111111101010","000000000000100000","111111111111111001","000000000000100001","000000000000001000","111111111111101000","111111111111101111","000000000000001101","000000000000010001","111111111111011110","000000000000001010","111111111111111100","111111111111110101","000000000000000011","111111111111010100","000000000000100101","111111111111110110","111111111111100000","000000000000010111","000000000000000011","000000000000000001","000000000000010010","000000000000101011","111111111111110000","111111111111110011","000000000000001100","000000000000000111","111111111111110011","000000000000010001","111111111111110000","000000000000000000","000000000000001101","000000000000001010","111111111111110101","111111111111111010","111111111111110010","111111111111111000","000000000000001110","111111111111101111","111111111111101100","000000000000001101","000000000000000000","000000000000001000","000000000000011100","111111111111110010","000000000000000001","111111111111100011","000000000000100100","000000000000001111","111111111111111001","000000000000000100","111111111111101010","000000000000100110","000000000000011010","111111111111011111","111111111111110010","111111111111111111","111111111110111101","000000000000011101","111111111111101001","111111111111010010","111111111111101010","111111111111101110","111111111111111010","111111111111101110","111111111111011001","111111111111110100","111111111111111010","111111111111111111","000000000000101001","000000000000000100","111111111111111100","111111111111101110","000000000000001111","000000000000001100","111111111111011101","000000000000010001","111111111111010010","111111111111110001","111111111111010100","000000000000001111","111111111111111110","111111111111011010","000000000000001110","000000000000010001","000000000000101101","111111111111011111","111111111111101111","111111111111110110","111111111111100110","111111111111101111","111111111111100110","000000000000000000","111111111111100110","111111111111011011","000000000000000000","111111111111110001","000000000000010001","111111111111111111"),
("000000000000010001","000000000000001010","111111111111011111","111111111111100010","111111111111110011","000000000000011001","111111111111111110","111111111111010010","111111111111111001","111111111111011111","111111111111001011","111111111111101110","000000000000010011","111111111111010010","000000000000000011","000000000000001011","111111111111111001","000000000000010111","111111111111110010","111111111111110111","000000000000001000","111111111111111100","000000000000001001","111111111111111000","000000000000010011","000000000000000001","111111111111011110","000000000000001100","111111111111111110","111111111111110010","000000000000010110","111111111111111001","000000000000010010","111111111111101011","111111111111110011","111111111111110011","111111111111111111","000000000000100100","111111111111001110","000000000000000000","111111111111111110","111111111111110100","111111111111101101","111111111110111000","000000000000101111","000000000000000010","111111111111100110","000000000000101001","000000000000011101","111111111111100101","000000000000010011","000000000000011101","000000000000000000","111111111111110011","000000000000010111","000000000000000101","111111111111110011","000000000000001000","111111111111110010","000000000000000000","111111111111111100","000000000000000101","111111111111111000","111111111111100011","111111111111100011","000000000000000011","000000000000011001","111111111111100101","111111111111100100","111111111111100111","000000000000001010","111111111111100001","000000000000010100","111111111111101101","000000000000000000","111111111111011111","000000000000100001","111111111111111010","111111111111110001","111111111111111001","000000000000000001","000000000000111111","000000000000001001","111111111111001010","111111111111111100","111111111111011100","111111111110010110","000000000000000101","111111111111101110","111111111111100100","000000000000000000","000000000000000111","000000000000000010","000000000000000001","111111111111001111","111111111111101110","111111111111111011","000000000000001101","000000000000111011","111111111111101100","000000000000001000","000000000000000101","111111111111111011","111111111111101111","111111111111110110","000000000000000100","111111111111110101","111111111111101100","111111111110111111","111111111111110111","000000000000001000","111111111111100001","000000000000000101","111111111111111110","000000000000000111","000000000000001101","000000000000001001","111111111111111011","111111111111010010","111111111111011101","000000000000001010","000000000000000111","111111111111100011","111111111110101110","111111111111111010","111111111111110111","111111111111110001","111111111111110001"),
("000000000000001010","000000000000101011","000000000000000111","111111111111111011","111111111111110100","000000000000001110","000000000000001101","111111111110110101","111111111111110101","111111111111111010","111111111111101100","111111111111001010","000000000000011100","111111111111111011","000000000000001101","000000000000001000","111111111111110111","000000000000010111","111111111111101000","111111111111111000","111111111111111000","000000000000000000","000000000000100000","000000000000001001","000000000000000111","000000000000000000","111111111111011000","111111111111111101","000000000000011001","111111111111110110","000000000000101001","111111111111100101","000000000000011011","111111111111111001","111111111111100101","111111111111111101","000000000000100001","000000000000010011","111111111111001101","000000000000000000","111111111111101100","111111111111101000","111111111111001010","111111111110111011","000000000000000010","111111111111110011","111111111111011000","000000000000010001","000000000000001000","111111111111110101","000000000000000111","000000000000000100","111111111111111101","111111111111100101","000000000000000000","000000000000000110","111111111111111001","000000000000001011","111111111111101111","111111111111111001","000000000000011000","000000000000011001","000000000000000101","000000000000000100","111111111111011110","000000000000000001","000000000000101100","000000000000001010","111111111111111011","111111111111110111","111111111111110101","111111111111110110","000000000000100001","111111111111101011","111111111111111011","111111111111101101","000000000000101001","111111111111111010","111111111111111101","000000000000010010","111111111111101111","000000000000100000","000000000000101010","111111111111111001","111111111111110111","111111111111101000","111111111110111100","000000000000000000","111111111111101001","111111111111011111","000000000000001111","000000000000001010","111111111111101100","111111111111110011","111111111111101011","111111111111001010","111111111111111101","000000000000100011","000000000000011010","000000000000000101","000000000000010010","111111111111000001","111111111111111001","000000000000000110","000000000000000000","000000000000000100","111111111111111001","111111111111011101","111111111110100110","000000000000010111","000000000000000111","000000000000000010","000000000000001111","000000000000000100","111111111111110011","000000000000010010","000000000000000001","111111111111101011","111111111111010100","111111111111110111","000000000000000110","000000000000011110","111111111111011000","111111111110101100","111111111111111101","000000000000001000","000000000000010101","111111111111110001"),
("000000000000011100","000000000000110011","111111111111110100","000000000000000011","111111111111101101","111111111111110111","000000000000100000","111111111111010110","111111111111111111","000000000000010010","111111111111110110","111111111111011000","000000000000010110","000000000000011100","111111111111101111","000000000000010011","000000000000011110","000000000000001100","111111111111110010","000000000000001111","111111111111110010","000000000000010000","000000000000011011","111111111111110011","111111111111111101","000000000000010111","111111111111101011","111111111111110000","111111111111110011","111111111111100010","000000000000011001","111111111111101111","000000000000000110","000000000000000000","111111111111111100","111111111111101011","111111111111111001","000000000000001001","111111111111000110","111111111111110111","111111111111000111","111111111111111000","111111111111000010","111111111111011010","000000000000001000","111111111111101111","111111111111100100","000000000000000011","000000000000000100","000000000000000011","000000000000010011","111111111111110101","000000000000001011","111111111111011100","000000000000001101","111111111111101100","000000000000000001","111111111111110011","000000000000011100","000000000000000011","000000000000001101","000000000000011110","000000000000001001","111111111111111010","111111111111101101","000000000000011010","000000000000000001","111111111111110110","111111111111100100","111111111111111100","000000000000010011","000000000000000111","000000000000100110","000000000000000110","111111111111100111","111111111111010111","000000000000000000","000000000000000000","000000000000001111","000000000000010110","111111111111110101","111111111111110001","000000000000010101","111111111111111111","111111111111101011","000000000000000101","111111111110010101","111111111111100010","111111111111110111","111111111111011111","000000000000011000","000000000000000110","111111111111111101","000000000000000110","111111111111010101","111111111111010010","000000000000001111","000000000000001000","000000000000011111","111111111111101101","000000000000000001","111111111111011100","111111111111111001","000000000000001001","000000000000010000","000000000000010100","111111111111110111","111111111111011101","111111111110111110","111111111111111001","000000000000001101","111111111111111000","111111111111111000","000000000000000111","111111111111100110","000000000000100000","000000000000000001","111111111111101001","111111111111001110","111111111111001110","111111111111111000","000000000000011001","111111111111010100","111111111110110110","000000000000000101","111111111111110111","000000000000000001","111111111111100000"),
("000000000000100010","000000000000100111","111111111111110010","111111111111111110","111111111111110110","000000000000011000","000000000000001111","111111111111100110","000000000000010011","000000000000001010","000000000000000111","111111111111011100","000000000000001110","000000000000011011","111111111111011000","000000000000000011","000000000000000101","000000000000000111","000000000000001001","000000000000000001","000000000000000011","000000000000010010","000000000000000000","000000000000100111","000000000000000001","000000000000011101","111111111111101111","111111111111111100","111111111111110100","111111111111001101","000000000000010010","111111111111111001","111111111111110011","111111111111101110","000000000000000111","111111111111111011","111111111111101100","000000000000010000","111111111111110101","111111111111100101","111111111111010111","111111111111111011","111111111111011010","000000000000001011","111111111111111100","111111111111110010","000000000000001100","111111111111101010","000000000000000000","111111111111111000","000000000000101101","111111111111111010","000000000000010001","111111111111100101","111111111111101000","111111111111110001","111111111111100010","111111111111101111","000000000000010110","111111111111101110","111111111111111101","000000000000010011","000000000000000110","000000000000011000","111111111111101001","000000000000001110","111111111111111110","000000000000000100","111111111111111101","111111111111110110","000000000000000111","111111111111110011","000000000000010000","111111111111101011","111111111111110000","111111111111010001","000000000000001111","111111111111111000","111111111111111111","111111111111111011","111111111111111110","111111111111100001","000000000000001011","000000000000010010","111111111111101011","111111111111111000","111111111110100011","111111111111100101","000000000000001010","111111111111110000","111111111111110001","111111111111101100","111111111111101111","000000000000010110","111111111111111000","111111111111001100","111111111111110100","111111111111101111","000000000000001000","111111111111110000","000000000000100100","111111111111111001","000000000000001110","000000000000000010","000000000000010101","000000000000001011","111111111111100100","111111111111101001","111111111111001111","000000000000000010","000000000000001000","111111111111111001","000000000000000001","000000000000000010","111111111111111110","000000000000100111","111111111111111001","111111111111010001","111111111111010101","111111111111000010","000000000000000110","000000000000011001","111111111111100101","111111111101111100","111111111111111110","111111111111110010","000000000000010110","111111111111111101"),
("000000000000100101","000000000000110000","111111111111110101","000000000000000000","111111111111110110","111111111111111110","000000000000001111","111111111111110100","000000000000001100","111111111111111010","000000000000100010","111111111111110001","000000000000001001","000000000000101011","111111111110111110","111111111111111101","000000000000001101","000000000000010001","000000000000101011","000000000000000101","000000000000001101","111111111111111011","000000000000011011","111111111111111110","111111111111101101","000000000000000110","000000000000100100","000000000000001101","111111111111011001","111111111111011101","000000000000011100","111111111111110101","000000000000000000","111111111111100100","000000000000000100","111111111111001000","111111111111110111","111111111111110011","111111111111101010","000000000000001011","111111111111010011","000000000000000101","000000000000011010","000000000000101100","000000000000011010","111111111111100001","000000000000111100","111111111111100011","111111111111110111","111111111111111100","000000000000001010","111111111111110011","000000000000010101","111111111111110001","111111111111110010","000000000000001010","111111111111100111","111111111111111000","000000000000000110","111111111111110100","111111111111110111","000000000000011011","000000000000000110","000000000000001101","111111111111001100","000000000000001001","000000000000011100","000000000000011000","111111111111111101","111111111111100000","000000000000010111","000000000000001101","000000000000011100","000000000000001110","111111111111010110","111111111111010011","000000000000011111","111111111111111100","111111111111100111","111111111111111100","111111111111110100","000000000000010111","000000000000000111","111111111111111111","111111111111110001","111111111111111001","111111111110010110","111111111111100001","000000000000001011","111111111111110110","111111111111101010","111111111111111101","000000000000010000","000000000000000010","000000000000010011","111111111111100101","111111111111110110","111111111111110010","111111111111110101","111111111111110010","000000000000001010","000000000000000000","000000000000010000","000000000000000000","000000000000001100","000000000000100100","111111111111100000","111111111111111011","111111111111100000","111111111111101110","111111111111101011","111111111111111000","000000000000000110","111111111111100001","000000000000011000","000000000000001001","000000000000000110","111111111111010111","111111111111011011","111111111111011110","000000000000000000","000000000000010001","111111111111101100","111111111110010000","000000000000010011","000000000000000100","000000000000001101","111111111111101100"),
("000000000000011001","000000000000001001","111111111111100100","000000000000001011","000000000000010000","111111111111111110","111111111111100000","000000000000011111","111111111111100110","000000000000000001","000000000000101010","000000000000000010","000000000000011010","000000000000110011","111111111111010111","000000000000000100","000000000000000000","000000000000000000","000000000000010100","000000000000000101","000000000000010110","000000000000000000","000000000000001001","000000000000010001","000000000000000010","000000000000001001","000000000000010010","000000000000001111","111111111111110111","111111111111100111","000000000000000110","000000000000000111","111111111111111011","111111111111111011","000000000000001001","111111111111100000","000000000000000111","000000000000001001","000000000000001101","111111111111111010","111111111111011000","000000000000010111","000000000000100001","000000000000010010","000000000000001110","111111111111010100","000000000000101010","111111111111001101","000000000000000100","111111111111100110","111111111111111100","000000000000000000","111111111111111101","111111111111010110","111111111111101000","111111111111111001","000000000000000000","000000000000010010","000000000000010011","111111111111110000","111111111111100101","000000000000001111","000000000000000000","000000000000001100","111111111111101101","000000000000001000","000000000000000010","000000000000001100","111111111111111111","111111111111110101","000000000000010000","111111111111110100","000000000000000000","111111111111101011","111111111111100101","111111111111010000","000000000000100001","111111111111111100","111111111111011011","000000000000001111","111111111111111100","000000000000010100","111111111111101100","000000000000000001","111111111111100011","000000000000001000","111111111110111101","111111111111100101","000000000000010001","111111111111110010","111111111111011001","111111111111100101","000000000000001001","111111111111101001","000000000000101010","111111111111110001","111111111111100011","000000000000010111","000000000000001010","000000000000001011","000000000000001011","111111111111111101","111111111111011001","000000000000000000","000000000000001010","000000000000010111","111111111111101111","000000000000101111","111111111111011000","111111111111101111","111111111111111011","111111111111111001","000000000000000010","111111111111101101","000000000000010110","000000000000010010","000000000000011000","111111111111011110","111111111111110110","111111111111011101","111111111111101101","000000000000011010","000000000000011000","111111111110011001","000000000000000010","000000000000000010","111111111111110001","000000000000000011"),
("000000000000010101","000000000000001111","111111111111100010","111111111111110100","111111111111110101","111111111111111101","111111111111110101","000000000000000100","000000000000000000","111111111111110001","000000000000110110","000000000000000111","000000000000001000","000000000000011000","111111111111010110","000000000000000100","111111111111111001","111111111111101011","000000000000101111","000000000000000100","111111111111110100","000000000000000010","000000000000001101","111111111111111110","111111111111101000","000000000000001110","000000000000101010","111111111111111010","000000000000001010","111111111111110101","000000000000001011","000000000000000000","111111111111110011","111111111111100101","000000000000101100","111111111111100001","111111111111111011","000000000000010000","000000000000010011","111111111111110010","111111111110111011","000000000000011001","000000000000111110","000000000000000000","000000000000101100","000000000000000111","000000000000100111","000000000000001110","111111111111110110","111111111111110011","111111111111010001","111111111111111011","111111111111100001","111111111110111100","111111111111100001","000000000000000011","000000000000000000","000000000000000100","111111111111101010","111111111111110101","111111111111101100","000000000000000011","111111111111111111","000000000000011011","111111111111110010","000000000000000000","000000000000000000","000000000000000000","000000000000000011","111111111111101001","000000000000010110","111111111111110010","000000000000001110","111111111111011110","111111111111001011","111111111111000101","000000000000010011","000000000000000010","111111111111111110","000000000000000111","000000000000000111","000000000000010100","000000000000001111","000000000000100100","111111111111100010","111111111111110100","111111111101111000","111111111111111101","000000000000110110","111111111111111111","111111111111001100","111111111111010011","111111111111111110","000000000000010010","000000000000001100","111111111111011001","111111111111011101","000000000000010100","000000000000100000","000000000000011011","000000000000000000","000000000000100111","111111111111110101","111111111111111111","000000000000000000","000000000000000101","111111111111110101","000000000000011110","111111111111101101","111111111111100100","111111111111100100","111111111111110001","000000000000100111","111111111111101110","000000000000000110","111111111111100111","000000000000011001","111111111111011001","111111111111101000","111111111111011101","000000000000001111","000000000000001101","000000000000100110","111111111111101001","111111111111111110","000000000000010101","000000000000000110","111111111111110001"),
("000000000000100001","111111111111111011","111111111111101111","000000000000001010","000000000000010011","000000000000100000","000000000000000101","000000000000010001","111111111111101101","111111111111101100","000000000000100000","000000000000000001","000000000000010010","000000000000111000","111111111111100111","111111111111111011","000000000000010011","111111111111111110","000000000000001100","111111111111110101","111111111111111000","111111111111010000","111111111111101011","000000000000010001","111111111111101001","000000000000011100","000000000000000000","000000000000001001","000000000000011111","111111111111100010","000000000000001010","111111111111111010","111111111111101010","111111111111101111","000000000000010110","111111111111100111","111111111111110110","000000000000010101","000000000000010100","111111111111110010","111111111110110000","000000000000100110","000000000000001010","000000000000001110","000000000000010000","000000000000000111","000000000000100011","000000000000000111","111111111111111000","111111111111110101","111111111111000110","000000000000001100","111111111111111010","111111111111001001","111111111111110010","000000000000011010","000000000000001001","111111111111111000","000000000000001010","111111111111111010","111111111111101011","000000000000000000","111111111111111000","000000000000000001","111111111111110100","111111111111101111","000000000000000011","000000000000001100","000000000000000110","000000000000000101","000000000000001011","000000000000001001","000000000000001011","111111111111110000","111111111111111001","111111111111011011","000000000000010110","111111111111110111","000000000000001000","000000000000001000","000000000000001101","000000000000000000","000000000000001100","000000000000000011","111111111111101000","111111111111111011","111111111101111011","000000000000000111","000000000000100111","000000000000000001","111111111111110000","111111111111011001","000000000000010010","000000000000011000","000000000000010100","111111111111010010","111111111111100110","000000000000000110","000000000000101001","000000000000000100","000000000000000110","000000000000101100","111111111111101000","111111111111101000","000000000000010010","000000000000001010","000000000000000101","000000000000010111","000000000000000000","111111111111111100","000000000000010010","111111111111101000","000000000000000101","000000000000000011","000000000000010011","111111111111111110","111111111111111101","111111111111101010","000000000000000010","111111111111011000","000000000000000011","111111111111101111","000000000000011111","000000000000100111","000000000000010101","111111111111101100","111111111111100100","000000000000010001"),
("000000000000000000","111111111111111011","000000000000000100","111111111111101100","111111111111101101","000000000000011111","000000000000000101","000000000000010000","111111111111111010","111111111111011110","000000000000001100","111111111111100111","000000000000011111","000000000000010010","000000000000001100","111111111111111101","000000000000011010","111111111111110110","111111111111110110","000000000000010000","111111111111111000","111111111111000100","000000000000000011","111111111111011110","111111111111110111","000000000000010011","111111111111100101","111111111111101110","000000000000001001","111111111111100001","000000000000011000","000000000000000111","111111111111100001","000000000000001010","000000000000001101","111111111111011100","000000000000011001","111111111111111101","000000000000001010","000000000000001010","000000000000000100","111111111111111010","000000000000000010","000000000000000011","111111111111111101","000000000000100011","000000000000010110","000000000000010011","000000000000001001","000000000000000010","111111111111101100","111111111111111011","111111111111110010","111111111111110001","111111111111111000","000000000000001000","000000000000100001","111111111111110000","000000000000000110","000000000000000111","111111111111111001","000000000000000000","000000000000000001","111111111111110100","000000000000001011","000000000000000000","000000000000011010","000000000000000001","111111111111100011","000000000000010100","000000000000000010","111111111111101011","000000000000110001","111111111111101111","111111111111110100","111111111111101111","000000000000010010","000000000000001010","000000000000001000","000000000000000011","111111111111111100","000000000000000101","000000000000011011","000000000000001010","111111111111101011","000000000000001110","111111111111000100","111111111111110001","111111111111101110","111111111111101100","000000000000011110","111111111111001000","000000000000001111","111111111111110111","111111111111101110","111111111111110000","111111111111010100","000000000000000101","000000000000000001","000000000000000101","111111111111110101","000000000000001010","111111111111100101","111111111111100110","111111111111100010","111111111111101111","000000000000001010","111111111111111001","111111111111110111","000000000000011001","000000000000001000","111111111111011101","111111111111111011","111111111111101101","000000000000000011","111111111111110111","000000000000000001","111111111111111100","000000000000010111","111111111111101000","111111111111110110","111111111111110110","000000000000000011","000000000001000110","000000000000010111","111111111111100001","111111111111101011","000000000000000000"),
("000000000000001110","111111111111011110","000000000000010011","000000000000000111","111111111111101110","111111111111111011","000000000000000000","111111111111111110","111111111111110000","111111111111111110","000000000000000010","111111111111001011","000000000000001010","111111111111100001","000000000000101011","000000000000000001","000000000000000010","000000000000000001","000000000000010011","000000000000010110","111111111111111000","111111111110110100","000000000000001010","111111111111110100","000000000000010001","000000000000001100","111111111111011111","111111111111110010","000000000000010110","111111111111101011","000000000000000100","000000000000001101","000000000000000110","000000000000001101","000000000000000011","111111111111100101","000000000000011010","000000000000100001","111111111111111110","000000000000011110","000000000000010101","111111111111111001","000000000000000000","111111111111100100","000000000000010101","000000000000000111","000000000000010010","000000000000010110","000000000000000111","000000000000001001","111111111111101111","000000000000001100","111111111111100101","000000000000011100","000000000000011000","000000000000001111","000000000000011000","000000000000001100","000000000000001001","111111111111110011","000000000000000011","111111111111110110","111111111111110000","111111111111110011","111111111111110110","111111111111111110","000000000000010000","000000000000001011","111111111111011110","111111111111101110","000000000000010001","000000000000001100","000000000000110001","000000000000000101","000000000000010000","000000000000010011","111111111111101101","000000000000000111","000000000000000000","000000000000001101","111111111111111000","111111111111101000","000000000000111110","111111111111111010","111111111111111111","000000000000010001","111111111111101000","111111111111111111","000000000000000000","000000000000000110","000000000000101101","111111111111101110","111111111111100001","111111111111110100","000000000000001011","000000000000001000","111111111111100101","111111111111110101","000000000000010000","111111111111111110","000000000000000100","000000000000010001","000000000000000110","000000000000000010","111111111111010100","111111111111111010","000000000000000010","000000000000001111","000000000000001001","000000000000011000","111111111111101111","111111111111101101","111111111111111100","000000000000010011","111111111111111111","000000000000000101","111111111111110010","000000000000000011","111111111111111001","111111111111111110","111111111111100111","111111111111111101","000000000000000001","000000000000111000","000000000000110000","111111111111101100","111111111111111000","000000000000011000"),
("111111111111111100","111111111111100100","000000000000010011","000000000000000110","111111111111101111","000000000000010101","111111111111110100","111111111111111001","111111111111101101","000000000000001100","000000000000001001","111111111111001001","000000000000001100","111111111111101001","000000000000100011","000000000000001100","000000000000100111","111111111111111010","111111111111111110","000000000000001010","111111111111110001","111111111111010111","000000000000100100","111111111111010111","111111111111111010","000000000000001010","111111111111111101","000000000000001101","000000000000001011","000000000000011001","000000000000000001","000000000000000100","000000000000011000","000000000000000011","111111111111101010","111111111111110101","111111111111111111","000000000000010110","000000000000000001","000000000000011101","000000000000010010","111111111111101001","111111111111111100","111111111111110001","000000000000011001","111111111111101101","000000000000011000","111111111111111111","111111111111111110","000000000000001111","111111111111101101","000000000000000101","111111111111110011","000000000000000001","111111111111111001","111111111111110011","000000000000001100","111111111111110111","000000000000000000","000000000000001010","000000000000001101","000000000000000011","111111111111110101","111111111111111101","111111111111010010","000000000000000000","000000000000101100","000000000000010001","000000000000000100","111111111111110000","111111111111101111","000000000000001100","000000000000011110","111111111111101111","111111111111110011","000000000000100100","000000000000001101","000000000000001011","111111111111111001","000000000000001100","111111111111110100","000000000000010101","000000000000100110","111111111111011111","111111111111110110","000000000000011000","000000000000100001","111111111111111101","111111111111110101","111111111111110101","000000000000001011","000000000000000000","000000000000000001","111111111111011100","000000000000001111","000000000000000111","111111111111111111","111111111111101111","111111111111111011","111111111111110110","111111111111111010","000000000000001010","000000000000011111","111111111111111111","111111111111110111","111111111111111101","000000000000001100","000000000000010100","000000000000010100","000000000000100100","000000000000000111","111111111111110111","000000000000011101","000000000000001010","000000000000001101","111111111111111000","000000000000001011","000000000000000111","000000000000010000","000000000000000100","111111111111111111","000000000000001110","111111111111101000","000000000000101101","000000000000111101","111111111111110110","000000000000001000","000000000000000011"),
("111111111111101100","000000000000000110","111111111111110100","111111111111111010","111111111111110000","000000000000001010","000000000000001001","111111111111101110","111111111111110110","000000000000000011","111111111111110100","111111111111101101","000000000000010001","111111111111100110","000000000000011110","111111111111111111","000000000000000111","000000000000001010","000000000000011101","000000000000000001","000000000000000100","000000000000000000","000000000000001010","111111111111100010","000000000000000011","111111111111111110","111111111111111001","111111111111111110","111111111111111110","000000000000001010","000000000000001001","000000000000010111","000000000000100010","000000000000001110","111111111111100110","111111111111110100","000000000000010100","000000000000010101","111111111111111011","111111111111111100","000000000000011001","111111111111101000","000000000000011001","111111111111110110","000000000000000010","111111111111101010","000000000000010100","000000000000101000","111111111111111011","111111111111111001","111111111111011011","111111111111110101","111111111111110111","000000000000011111","111111111111111000","111111111111101101","000000000000010111","000000000000001111","111111111111111111","000000000000001101","000000000000001000","111111111111100100","000000000000001101","111111111111101010","111111111110101101","000000000000001101","000000000000000011","000000000000000011","000000000000010001","111111111111110000","111111111111111111","111111111111111111","000000000000100101","000000000000001110","000000000000010110","000000000000100100","111111111111111010","111111111111101010","000000000000000110","111111111111111100","000000000000010000","111111111111111001","000000000000011100","000000000000000011","000000000000000000","000000000000001000","000000000000100100","000000000000001000","000000000000000100","000000000000010010","000000000000010101","000000000000010101","111111111111111010","111111111111110010","000000000000000100","000000000000010110","000000000000000100","000000000000001001","000000000000000110","111111111111101011","111111111111111100","111111111111100110","000000000000101000","111111111111110110","111111111111101000","111111111111100111","111111111111100100","000000000000010110","111111111111110101","000000000000000000","111111111111101011","000000000000001110","000000000000000011","111111111111111000","111111111111111011","000000000000000010","000000000000011010","111111111111111100","111111111111111101","000000000000001100","111111111111100110","000000000000001011","111111111111010100","000000000000011001","000000000000101010","111111111111110000","111111111111111011","000000000000001100"),
("111111111111101110","000000000000010010","111111111111101001","111111111111110011","111111111111110010","111111111111110100","000000000000000110","000000000000000110","111111111111111010","000000000000010111","111111111111110101","111111111111111010","111111111111110101","111111111111010100","000000000000000101","111111111111111111","000000000000000111","111111111111111011","111111111111110111","111111111111111110","111111111111111111","000000000000010010","000000000000110011","111111111111111011","111111111111111001","000000000000010100","000000000000000000","111111111111111010","000000000000010011","000000000000101011","111111111111101111","000000000000001010","000000000000011000","000000000000000011","111111111111101001","111111111111111110","000000000000010001","111111111111111110","000000000000001010","000000000000000101","111111111111110111","111111111111110110","000000000000011000","111111111111110001","000000000000000110","111111111111100100","000000000000101010","000000000000001100","000000000000001000","000000000000001100","111111111111011101","111111111111110111","111111111111111110","000000000000000001","000000000000001000","111111111111101100","000000000000010000","111111111111110111","000000000000000110","111111111111110101","111111111111111110","111111111111100111","000000000000011100","111111111111111101","111111111110110011","111111111111111010","111111111111110010","111111111111110101","000000000000001000","000000000000001101","000000000000001000","111111111111110000","000000000000011010","000000000000000011","000000000000010011","000000000000000110","000000000000010000","111111111111100000","000000000000000011","000000000000000011","000000000000001011","000000000000011001","000000000000101100","111111111111111100","111111111111110111","000000000000000100","000000000000000101","000000000000000111","000000000000001001","000000000000000011","000000000000010000","000000000000010011","111111111111101100","000000000000011000","000000000000001100","000000000000010100","111111111111111010","000000000000010100","000000000000010100","000000000000000101","111111111111111100","111111111111111011","000000000000001001","111111111111110100","000000000000001000","111111111111110000","111111111111110111","111111111111110100","111111111111110100","000000000000000000","111111111111110101","000000000000010110","111111111111111000","111111111111111010","111111111111111010","000000000000000111","111111111111110011","000000000000000111","111111111111101011","000000000000001011","000000000000000010","111111111111111011","111111111111110001","000000000000100011","000000000000100011","111111111111110111","111111111111111001","111111111111111100"),
("111111111111110001","000000000000110001","111111111111101100","111111111111110011","111111111111100011","111111111111111110","111111111111100100","000000000000110111","000000000000000000","000000000000001100","111111111111111100","000000000000010001","111111111111110101","111111111111101011","111111111111111111","111111111111111100","111111111111110001","111111111111101110","000000000000000100","000000000000010010","111111111111111101","111111111111110010","000000000000000010","111111111111100011","000000000000001001","111111111111111100","111111111111110101","000000000000000100","000000000000010101","111111111111111101","111111111111111110","111111111111110111","000000000000010010","000000000000001010","111111111111101000","000000000000001100","000000000000000010","000000000000011001","000000000000001100","000000000000100011","000000000000001111","111111111111101001","000000000000001100","111111111111100101","000000000000010111","111111111111100010","000000000000000110","000000000000000100","000000000000011101","111111111111101001","111111111111001011","000000000000000101","111111111111100101","000000000000100110","111111111111111111","111111111111111110","000000000000001011","111111111111110100","000000000000001101","111111111111101110","000000000000011110","111111111111111101","000000000000011111","111111111111111011","111111111111001011","000000000000000101","111111111110111000","111111111111111011","000000000000010010","111111111111101110","111111111111111110","000000000000001101","111111111111111111","111111111111111100","000000000000010101","000000000000101000","111111111111110010","000000000000000100","000000000000001001","111111111111101000","111111111111100010","000000000000100010","000000000000001000","000000000000001000","111111111111110101","000000000000000000","000000000000000110","000000000000001111","111111111111110101","000000000000010110","111111111111111001","000000000000100110","111111111111111010","000000000000000010","111111111111101010","111111111111101011","111111111111111010","111111111111110101","000000000000010101","111111111111101101","111111111111110101","111111111111101000","111111111111111110","111111111111111011","111111111111110011","111111111111101010","111111111111111110","111111111111101101","111111111111101000","000000000000001010","111111111111111000","111111111111111000","000000000000001111","111111111111110101","111111111111101111","111111111111110000","000000000000010011","111111111111101011","111111111111110000","000000000000011000","111111111111110010","000000000000000101","111111111111011011","000000000000011000","000000000000011001","000000000000000111","111111111111100000","000000000000000000"),
("111111111111110101","000000000000011011","111111111111101110","111111111111011011","000000000000000110","000000000000010010","111111111111101111","000000000000010010","000000000000000011","111111111111111101","111111111111110100","000000000000011011","111111111111111000","000000000000000010","000000000000000101","111111111111111011","111111111111110011","111111111111110010","111111111111110100","000000000000010001","000000000000000000","111111111111111010","111111111111111000","111111111111101000","000000000000000101","111111111111111011","111111111111010011","111111111111110000","111111111111111101","111111111111011011","111111111111111001","111111111111110001","000000000000000011","000000000000011010","111111111111110111","000000000000000110","000000000000001000","000000000000000011","111111111111111000","000000000000001110","000000000000010011","000000000000000101","000000000000000000","111111111111100100","111111111111110011","111111111111111101","111111111111111110","000000000000001001","000000000000010001","000000000000001001","111111111111111010","000000000000001101","111111111111111101","000000000000010001","000000000000000011","000000000000000101","111111111111110100","111111111111110001","000000000000010001","111111111111101111","111111111111111010","000000000000000000","000000000000001010","111111111111110011","111111111111000100","000000000000001100","111111111110110111","111111111111111000","000000000000010110","000000000000010110","111111111111110001","000000000000000011","111111111111010110","000000000000011010","000000000000011001","000000000000100001","000000000000010010","111111111111110110","111111111111110011","000000000000000000","111111111111110111","000000000000001110","000000000000011000","111111111111100100","000000000000001011","111111111111101100","000000000000001000","000000000000011000","000000000000000110","000000000000010101","111111111111111011","111111111111110010","111111111111111000","000000000000011000","111111111111101100","111111111110111101","111111111111111010","111111111111111001","111111111111110000","111111111111111101","000000000000010101","000000000000001000","111111111111010110","000000000000001111","000000000000000000","111111111111111001","000000000000000101","111111111111101000","111111111111011011","111111111111110000","000000000000010010","000000000000000011","000000000000010110","111111111111110100","000000000000000000","111111111111111000","111111111111101001","000000000000000000","111111111111001000","111111111111111111","111111111111111110","000000000000000100","000000000000001001","000000000000000110","111111111111111010","000000000000000000","000000000000000011","000000000000000110"),
("000000000000001011","000000000000100001","111111111111101100","111111111111111100","000000000000011010","000000000000001010","111111111111110001","000000000000100011","111111111111100000","000000000000000010","111111111111111100","000000000000001111","111111111111011110","111111111111101100","111111111111110101","111111111111110111","000000000000000100","000000000000000011","111111111111110010","111111111111111111","000000000000001000","111111111111111010","000000000000010110","111111111111101101","111111111111111100","111111111111101100","111111111111101110","111111111111110011","000000000000011010","111111111111110111","000000000000001010","111111111111110100","111111111111101011","000000000000000010","000000000000001100","111111111111110100","000000000000000111","000000000000000100","111111111111101110","000000000000010010","000000000000011111","000000000000011011","111111111111110101","111111111111101000","000000000000001101","000000000000010110","111111111111110101","000000000000010001","000000000000000000","111111111111101110","000000000000010100","000000000000000000","000000000000000011","000000000000010101","000000000000000111","000000000000001101","111111111111100011","000000000000000001","000000000000000001","111111111111111001","111111111111101111","111111111111110100","000000000000011111","111111111111110101","111111111111110001","111111111111101110","111111111110101010","111111111111111001","000000000000010100","111111111111101011","111111111111110110","111111111111111110","111111111110101010","000000000000011010","000000000000001000","000000000000100100","000000000000000011","111111111111101001","111111111111101100","000000000000010000","111111111111110111","000000000000000001","000000000000010100","111111111111000011","111111111111110101","111111111111111010","111111111111111000","000000000000011010","000000000000010101","000000000000001100","111111111111110011","111111111111110010","111111111111111011","000000000000001110","111111111111110101","111111111110111011","111111111111111101","000000000000010001","111111111111110010","111111111111111100","000000000000000000","111111111111011101","111111111111100000","111111111111101010","000000000000000000","000000000000001101","000000000000000000","111111111111101001","111111111111101110","111111111111111110","111111111111111011","111111111111100011","000000000000000001","000000000000010111","111111111111111000","111111111111100110","111111111111110001","000000000000100010","111111111111101011","000000000000011111","000000000000010100","000000000000001000","000000000000000111","111111111111110010","000000000000001110","111111111111110101","000000000000001000","111111111111111111"),
("000000000000000010","000000000000101100","111111111111110101","000000000000000100","111111111111110010","000000000000000100","111111111111111111","000000000000000011","111111111111101111","000000000000011001","000000000000000010","000000000000100111","111111111111111101","111111111111101011","111111111111101110","000000000000010100","000000000000000001","111111111111111100","111111111111111101","000000000000011011","000000000000010001","000000000000000000","000000000000011000","111111111111100011","111111111111101101","111111111111101100","111111111111101011","111111111111101010","111111111111110001","111111111111100011","111111111111110110","111111111111101000","000000000000001111","111111111111010010","111111111111111001","111111111111111011","000000000000001100","000000000000011010","111111111111100110","111111111111111001","000000000000001001","111111111111110101","111111111111110111","111111111111010110","111111111111101100","111111111111110010","000000000000000100","000000000000000101","111111111111110010","111111111111111111","000000000000011101","111111111111110001","000000000000001000","000000000000000100","000000000000011001","111111111111101101","111111111111000101","111111111111111100","000000000000001111","000000000000010001","111111111111100111","111111111111111011","000000000000011111","111111111111111110","000000000000000000","000000000000000011","111111111110111110","111111111111111010","111111111111111111","111111111111111111","000000000000011000","111111111111110011","111111111111001010","000000000000001011","000000000000001110","000000000000011111","111111111111101011","111111111111100100","111111111111110011","111111111111110110","111111111111011101","111111111111100010","000000000000001101","111111111110110111","000000000000010001","111111111111110101","000000000000000110","000000000000100110","000000000000000110","000000000000001110","111111111111101110","000000000000001100","000000000000001011","000000000000010000","111111111111111110","111111111111101101","000000000000000001","111111111111101100","111111111111100001","111111111111101111","000000000000010001","111111111111100110","111111111111101111","000000000000001111","111111111111110011","000000000000000110","000000000000000100","111111111111110110","111111111111011101","111111111111011000","111111111111111011","111111111111110100","111111111111110100","000000000000000101","000000000000000111","000000000000001000","111111111111111100","000000000000000000","111111111111001001","000000000000001100","111111111111111100","111111111111111111","000000000000010011","111111111111111100","000000000000010011","111111111111111000","111111111111111011","111111111111111000"),
("000000000000001111","000000000000000101","000000000000001100","111111111111101110","111111111111100010","000000000000011011","000000000000000111","111111111111101001","000000000000001010","111111111111110110","000000000000001101","000000000000100111","111111111111101001","000000000000000010","111111111111011111","111111111111111111","000000000000001110","111111111111110111","111111111111111110","111111111111111100","000000000000010101","111111111111110011","000000000000001010","111111111111111010","000000000000000100","000000000000010100","000000000000010110","000000000000010011","111111111111111001","111111111111100011","000000000000010001","111111111111100100","000000000000000101","111111111111001001","000000000000000001","000000000000001011","111111111111110001","000000000000010110","111111111111010010","111111111111111001","000000000000001111","111111111111111111","000000000000001100","111111111111111011","111111111111110111","111111111111101110","000000000000010110","000000000000100001","111111111111101101","111111111111110001","000000000000110001","111111111111110110","111111111111111001","111111111111110011","000000000000010001","111111111111100100","111111111111100100","000000000000000010","111111111111100010","000000000000000000","111111111111010011","111111111111110101","000000000000011001","000000000000000011","000000000000010101","111111111111100010","111111111111011000","111111111111111101","000000000000000000","111111111111110000","111111111111111011","000000000000000101","111111111111110001","111111111111100111","000000000000000011","000000000000001100","000000000000001111","111111111111100010","111111111111100110","000000000000000011","111111111111011101","111111111111110101","000000000000010101","111111111111000000","000000000000000010","111111111111000100","111111111111101100","000000000000011010","000000000000011010","111111111111101100","000000000000010000","111111111111111000","111111111111111100","111111111111110001","111111111111101000","111111111111001101","000000000000010000","000000000000000111","111111111111011001","111111111111011100","111111111111110110","111111111111111001","111111111111101010","000000000000000011","111111111111100110","000000000000011111","111111111111101110","111111111111111000","111111111111011100","111111111111111010","111111111111101101","111111111111100011","000000000000010001","000000000000011100","111111111111100100","000000000000011101","111111111111101010","000000000000000101","111111111111001100","000000000000000001","000000000000001000","000000000000000000","000000000000011011","111111111111110000","000000000000010011","000000000000000000","111111111111110011","111111111111101010"),
("000000000000000000","111111111111111111","111111111111101010","111111111111110111","111111111111111011","000000000000000010","000000000000001111","111111111111101010","000000000000001011","111111111111111000","000000000000011100","000000000000010011","000000000000011001","111111111111111001","111111111111101010","000000000000011111","111111111111110001","000000000000010010","111111111111100001","111111111111110000","111111111111111110","111111111111100101","111111111111111101","111111111111111100","111111111111110001","111111111111111111","000000000000011101","000000000000001101","000000000000000001","111111111111010011","000000000000000011","111111111111110101","111111111111110011","111111111111011001","000000000000011111","111111111111101110","000000000000001000","000000000000011001","111111111111100110","111111111111111000","000000000000000111","111111111111110011","000000000000001100","000000000000000100","111111111111111100","111111111111100010","111111111111011011","000000000000100100","000000000000000000","111111111111101100","000000000000000111","000000000000000010","000000000000000000","000000000000000111","000000000000100111","111111111111110010","111111111111101100","111111111111111101","111111111111011110","111111111111110111","111111111111011001","000000000000001101","000000000000001111","111111111111101000","000000000000000000","111111111111100001","111111111111110110","111111111111011101","111111111111101100","111111111111101101","111111111111101110","111111111111110011","111111111111100101","111111111111101010","111111111111111100","000000000000000000","000000000000010000","111111111111110011","111111111111100011","111111111111101011","111111111111110111","111111111111110110","000000000000001111","111111111110111011","000000000000001110","111111111111010001","000000000000001011","000000000000001000","111111111111100011","111111111111011100","000000000000100001","111111111111101111","111111111111111111","000000000000011000","000000000000000010","111111111111001011","000000000000000111","111111111111011110","111111111111010000","111111111111100110","000000000000010100","000000000000010000","111111111110110111","111111111111101100","111111111111111100","000000000000000000","111111111111011110","111111111111100011","111111111111011110","111111111111100011","111111111111111111","111111111111100111","111111111111101001","111111111111110100","111111111111010011","000000000000010000","111111111111101000","000000000000010000","111111111111011001","111111111111100110","000000000000001010","000000000000010010","000000000000011110","111111111111111011","000000000000101100","000000000000000000","000000000000001110","111111111111001010"),
("000000000000100000","111111111111101100","111111111111110000","000000000000000111","000000000000000001","000000000000110110","000000000000000000","000000000000000011","000000000000100111","111111111111101001","000000000000000011","111111111111011010","000000000000001110","111111111111111001","111111111111111100","000000000000101011","000000000000010000","000000000000011011","111111111111010011","000000000000000011","000000000000011100","111111111111101110","111111111111111101","111111111111110110","111111111111011111","000000000000110000","000000000000000000","000000000000001011","000000000000011100","111111111111110101","000000000000001111","111111111111111011","111111111111110000","111111111111010110","000000000000110010","111111111111001111","000000000000000101","000000000000001001","111111111111100101","111111111111011101","111111111111110010","111111111111101111","000000000000110010","000000000000111001","111111111111001111","111111111111010111","000000000000001100","000000000000100001","111111111111001111","111111111111100001","111111111111111011","111111111111011001","111111111111100101","000000000000010110","000000000000101011","111111111111110110","111111111111101001","111111111111111110","111111111111100001","000000000000000001","111111111111100100","000000000000001000","000000000000011010","111111111111101111","000000000000010111","111111111111001000","000000000000000000","000000000000001010","000000000000100100","000000000000010000","000000000000100110","111111111111110010","000000000000011000","000000000000000101","111111111111111111","111111111111111101","000000000000001011","000000000000011100","111111111111101110","111111111111110101","000000000000000000","111111111111111101","000000000000101101","111111111111011001","111111111111111110","111111111111100101","000000000000010100","000000000000000110","111111111111101011","111111111111110010","111111111111111001","111111111111001001","111111111111110111","000000000000101000","111111111111110110","000000000000001100","111111111111101100","000000000000001011","000000000000001000","000000000000011000","000000000000100000","111111111111100001","111111111111010101","111111111111010101","000000000000001100","000000000000000111","111111111111010011","000000000000000111","111111111111011000","111111111111100100","111111111111101100","000000000000010011","111111111111101110","111111111111001011","111111111111011101","000000000000110111","000000000000000011","000000000000100110","000000000000000011","111111111111111111","000000000000011010","000000000000100011","000000000000010010","111111111111110000","000000000000111100","000000000000000110","000000000000011010","111111111111110000"),
("000000000000000000","111111111111001000","111111111111111011","000000000000000010","000000000000010000","000000000000001011","111111111111110100","000000000000000111","000000000000011100","111111111111101100","000000000000000100","111111111111100111","000000000000101100","000000000000001101","111111111111110100","000000000000001011","111111111111111111","000000000000011110","000000000000010100","000000000000010010","000000000000001111","111111111111110111","111111111111100100","000000000000011011","111111111111011100","000000000000000011","111111111111111010","000000000000000100","000000000000101101","000000000000001101","000000000000011001","000000000000001001","000000000000000000","111111111111110110","000000000000101010","111111111111111010","000000000000011110","111111111111101100","111111111111111101","000000000000100011","111111111111011000","000000000000010000","000000000000100111","111111111111110111","111111111111010100","111111111111111110","000000000000001110","000000000000001010","000000000000000101","111111111111110110","111111111111100101","111111111111110101","111111111111101011","000000000000001010","000000000000100101","000000000000011100","000000000000000001","000000000000011011","000000000000001110","111111111111110011","111111111111101001","000000000000100010","000000000000100001","111111111111111100","000000000000100110","111111111111110011","000000000000010000","111111111111010111","000000000001000011","111111111111101010","111111111111111010","000000000000000100","000000000000000011","000000000000111010","111111111111100101","111111111111101010","000000000000000101","111111111111100110","000000000000001101","000000000000010001","111111111111110110","111111111111100101","111111111111111100","000000000000100110","111111111111101111","111111111111111011","111111111111110100","111111111111110100","111111111111101000","000000000000000000","111111111111101000","111111111111111001","111111111111111100","000000000000000110","000000000000010110","111111111111110110","111111111111100101","111111111111111110","111111111111110101","000000000000001000","111111111111110100","111111111111010001","111111111111101101","111111111111011110","000000000000011101","111111111111110000","000000000000010100","000000000000000010","000000000000001011","111111111111110001","000000000000011011","000000000000011101","111111111111011000","111111111111110110","000000000000010111","000000000000000111","111111111111110111","000000000000100011","000000000000100101","111111111111111000","000000000000100101","111111111111110101","000000000000000011","000000000000011111","000000000000001000","111111111111001001","000000000000010001","000000000000000110"),
("000000000000110011","111111111111001011","000000000000001101","000000000000000001","000000000000011010","000000000000011010","000000000000101001","000000000000111001","000000000000011101","111111111111101111","000000000000011000","111111111111011111","000000000000101101","000000000000000011","111111111111110111","000000000000010100","000000000000101101","000000000000011001","111111111111101110","000000000000011000","000000000000010011","000000000000001110","111111111111110110","111111111111101101","111111111111011111","000000000000110011","111111111111111010","000000000000011001","000000000000011100","111111111111101100","000000000000011100","000000000000000100","000000000000010101","111111111111010001","000000000000100010","000000000000001110","000000000000010011","000000000000100010","000000000000000111","000000000000000000","111111111111010011","000000000000000011","000000000000110000","000000000000010110","000000000000011100","111111111111111110","111111111111111010","000000000000000110","111111111111100101","111111111111111000","111111111111101001","000000000000101000","111111111111011111","000000000000100000","000000000000101111","000000000000000010","111111111111110101","111111111111111001","111111111111110000","000000000000000110","111111111111111000","000000000000011110","000000000000011001","000000000000011000","000000000000100010","111111111111101100","000000000000000000","111111111111110111","000000000000000100","111111111111110010","000000000000011001","000000000000011000","000000000000100010","000000000000011011","111111111111100011","000000000000010100","000000000000101011","111111111111110111","111111111111111111","000000000000011100","000000000000000110","000000000000000110","000000000000101110","000000000000011000","111111111111110111","000000000000011101","000000000000001000","000000000000100100","111111111111110101","111111111111111110","111111111111110101","111111111111110000","111111111111100100","111111111111111101","111111111111110111","111111111111110011","000000000000000011","000000000000000010","111111111111100111","111111111111101011","000000000000101111","111111111111110110","000000000000000000","111111111111100100","000000000000000111","000000000000100001","111111111111100001","000000000000000000","000000000000100101","111111111111110010","111111111111100010","000000000000011111","000000000000001110","111111111111110011","111111111111101101","000000000000011000","000000000000001011","000000000000100111","111111111111111011","000000000000100100","000000000000011110","000000000000011010","000000000000010111","111111111111110011","000000000000111110","111111111111101000","000000000000101100","000000000000010000"),
("000000000000000110","000000000000000000","111111111111110101","111111111111110010","111111111111111111","000000000000000011","111111111111101101","111111111111111100","111111111111110110","000000000000001110","000000000000000010","111111111111101100","111111111111111000","111111111111110011","111111111111101110","111111111111101110","111111111111110000","000000000000001000","000000000000000000","111111111111101111","000000000000010010","111111111111111000","000000000000000001","000000000000010001","000000000000001100","000000000000000101","000000000000010001","000000000000000011","000000000000000000","000000000000000111","111111111111111011","111111111111111101","000000000000000100","111111111111111100","000000000000000010","000000000000010000","000000000000000000","000000000000010110","000000000000000111","000000000000001110","000000000000001011","000000000000010010","111111111111110001","111111111111111101","000000000000001001","111111111111110100","111111111111111010","000000000000000100","111111111111111111","111111111111111001","000000000000000011","000000000000001101","000000000000001111","000000000000001111","111111111111101111","000000000000001001","111111111111111001","111111111111110100","000000000000001000","111111111111110000","000000000000000110","000000000000001101","000000000000001000","000000000000010101","111111111111110100","000000000000010000","111111111111110001","111111111111110000","000000000000000000","111111111111110101","111111111111110111","111111111111111001","000000000000010101","111111111111101111","000000000000000011","111111111111101110","000000000000000011","000000000000000000","000000000000010000","111111111111111111","000000000000010100","111111111111110000","000000000000001110","000000000000010111","000000000000010000","000000000000010000","111111111111111010","111111111111111001","000000000000001001","000000000000010100","111111111111110000","111111111111110110","000000000000000000","000000000000010000","111111111111110111","111111111111110000","111111111111110001","111111111111111111","111111111111111010","000000000000000000","111111111111110000","111111111111111101","111111111111110011","111111111111111011","111111111111101110","111111111111101111","111111111111110000","111111111111101011","000000000000001101","111111111111111001","000000000000000001","111111111111110111","111111111111110001","000000000000000101","000000000000000001","000000000000000010","111111111111110100","111111111111110111","111111111111110100","000000000000000010","000000000000010010","111111111111111001","111111111111110011","111111111111110001","000000000000000010","000000000000001111","000000000000001001","000000000000000110"),
("111111111111100001","111111111111111110","000000000000000000","000000000000010001","111111111111111100","111111111111100100","000000000000010101","000000000000010011","000000000000010101","000000000000010110","000000000000001110","111111111111101111","000000000000010011","000000000000000111","000000000000011110","000000000000001001","111111111111110000","000000000000001010","111111111111111100","000000000000001010","000000000000100010","111111111111111011","111111111111111010","000000000000000111","000000000000001001","111111111111110100","111111111111101011","000000000000010000","111111111111111000","111111111111111111","111111111111111110","000000000000100110","000000000000001111","000000000000001110","000000000000001001","111111111111111001","000000000000100101","111111111111011111","111111111111100100","000000000000010000","000000000000001101","000000000000001111","000000000000010010","000000000000000100","111111111111110100","000000000000010010","000000000000010101","111111111111111000","000000000000000011","000000000000100000","000000000000101101","111111111111110011","000000000000010010","000000000000010010","000000000000001111","111111111111111110","111111111111101110","000000000000010010","000000000000010001","000000000000001001","000000000000110001","000000000000011100","000000000000000000","111111111111100111","111111111111100010","000000000000000001","000000000000100010","111111111111110110","111111111111110101","000000000000010011","111111111111111000","000000000000000100","000000000000001011","000000000000010101","111111111111111100","111111111111111110","111111111111101011","111111111111110101","000000000000001111","000000000000000000","111111111111110010","111111111111101001","000000000000000100","000000000000000010","111111111111110001","000000000000010001","000000000000010110","111111111111111011","111111111111110001","000000000000010110","000000000000000100","111111111111101001","000000000000010100","000000000000010100","000000000000100101","000000000000000000","111111111111110111","000000000000001100","000000000000001110","000000000000010010","111111111111101110","111111111111011101","111111111111110100","111111111111011000","000000000000011110","111111111111111000","111111111111011100","000000000000000011","111111111111011111","111111111111110101","000000000000001100","000000000000000110","111111111111011001","111111111111111111","111111111111111111","000000000000000111","000000000000000000","000000000000010001","111111111111110100","000000000000011001","000000000000000001","000000000000001111","000000000000010011","000000000000110000","000000000000010000","000000000000000110","111111111111111001","111111111111101001"),
("111111111111101111","000000000000001010","000000000000000110","111111111111110111","000000000000000011","111111111111101110","111111111111100001","000000000000000111","111111111111100111","000000000000000011","111111111111110100","000000000000010101","111111111111100111","000000000000100100","000000000000001000","111111111111110110","000000000000000000","000000000000001111","000000000000000100","000000000000000001","000000000000001011","000000000000011110","111111111111110000","111111111111110011","111111111111110110","111111111111101010","111111111111011001","111111111111111010","000000000000000000","111111111111111110","000000000000010101","111111111111110010","111111111111111010","000000000000010111","000000000000010011","111111111111110101","000000000000010010","111111111111111011","000000000000010011","000000000000000011","000000000000101000","000000000000010010","111111111111011111","111111111111110011","000000000000001011","111111111111110010","000000000000000000","111111111111111000","000000000000000111","000000000000000000","111111111111111111","111111111111110001","000000000000000011","000000000000000101","000000000000000011","111111111111110101","000000000000010101","000000000000000111","111111111111100010","111111111111101101","111111111111110111","111111111111111110","111111111111100011","111111111111100011","111111111111010010","000000000000001011","111111111111111000","000000000000000001","111111111111111110","111111111111110110","111111111111010110","111111111111101110","111111111111101110","111111111111101100","111111111111111101","111111111111110111","000000000000000110","111111111111111111","111111111111111010","111111111111111011","000000000000000111","111111111111110111","111111111111110000","111111111111110011","111111111111100100","111111111111111010","000000000000101011","000000000000000101","000000000000001101","111111111111110111","000000000000001110","111111111111110111","000000000000010001","111111111111101001","111111111111100110","111111111111101110","111111111111110100","000000000000001010","111111111111111111","000000000000000100","111111111111110110","111111111111001000","111111111111101001","111111111111010110","000000000000001010","111111111111100110","111111111111111011","111111111111111101","111111111111111110","111111111111111110","000000000000001111","000000000000011011","111111111111011101","111111111111101100","000000000000000000","111111111111011100","111111111111101011","000000000000011101","111111111111110011","111111111111110100","000000000000001010","000000000000000101","111111111111111111","000000000000010110","000000000000001011","000000000000010110","111111111111110100","000000000000001010"),
("111111111111111110","000000000000100001","111111111111110001","111111111111101101","000000000000011001","111111111111111100","111111111111001111","111111111111111001","000000000000001111","111111111111101010","111111111111111000","111111111111111100","111111111111110111","111111111111100000","111111111111010001","111111111111100100","000000000000110001","111111111111110101","000000000000000100","000000000000000101","111111111111100101","111111111111000110","000000000000001101","111111111111011000","111111111111110101","000000000000000010","111111111111110001","000000000000001110","000000000000000010","111111111111110111","111111111111111100","111111111111111010","000000000000100001","000000000000010111","111111111111110111","000000000000001111","111111111111111100","000000000000010111","111111111111111011","000000000000100000","000000000000010000","111111111111111011","111111111111110010","111111111111101101","000000000000101000","000000000000010100","111111111111110110","000000000000000000","000000000000001010","000000000000010110","111111111111101100","000000000001000010","111111111111001111","111111111111110011","000000000000001100","000000000000011010","000000000000001001","111111111111101101","111111111111110001","000000000000010011","111111111111111010","000000000000011001","000000000000010011","111111111111110101","000000000000000111","111111111111011010","111111111110111001","000000000000000001","111111111111000101","111111111111111011","000000000000000010","000000000000000111","111111111111010101","111111111111101000","000000000000001111","000000000000011100","000000000000000000","000000000000001101","111111111111110100","000000000000100111","000000000000001011","000000000000011010","000000000000101100","000000000000001110","111111111111111110","000000000000001110","000000000000001110","000000000000100011","000000000000010110","111111111111111010","000000000000001110","000000000000010011","111111111111110010","111111111111011111","111111111111001101","000000000000001100","000000000000001011","000000000000000100","000000000000110001","000000000000000110","000000000000001000","111111111111011011","111111111111110101","111111111111011011","111111111111111000","111111111111111001","111111111111100100","111111111111001110","111111111111111010","111111111111110011","111111111111100010","111111111111111100","000000000000011110","000000000000010111","000000000000001010","000000000000000000","111111111111110100","000000000000101110","111111111111110010","000000000000101001","000000000000010000","111111111111111101","000000000000000000","111111111111000010","000000000000101000","000000000000000001","111111111111110110","000000000000001011"),
("111111111111111000","000000000000000101","111111111111000001","111111111111111100","111111111111110001","000000000000010001","111111111111100101","111111111111111111","111111111111111110","000000000000000111","111111111111101011","111111111111111100","000000000000001001","111111111111011111","111111111111110010","111111111111110101","000000000000101011","000000000000000010","000000000000010111","111111111111111101","111111111111111111","000000000000010001","111111111111110000","111111111111010110","111111111111111110","000000000000001010","111111111111110100","111111111111110111","000000000000010111","000000000000000001","000000000000011010","000000000000000010","000000000000011010","000000000000000111","111111111111101001","111111111111100100","000000000000010111","000000000000101111","111111111111110111","000000000000010010","000000000000000011","000000000000000111","111111111111111111","111111111111100110","000000000000011111","111111111111100111","111111111111101010","000000000000010101","000000000000010001","111111111111111000","000000000000000000","000000000000010100","000000000000000000","000000000000001110","000000000000000110","000000000000001001","111111111111111101","111111111111111011","000000000000000110","111111111111111100","111111111111101110","000000000000000000","000000000000010001","000000000000001111","000000000000001000","111111111111111011","111111111111111111","111111111111111011","111111111111100101","000000000000011001","111111111111110110","000000000000001010","000000000000001010","111111111111110111","000000000000001110","111111111111110011","000000000000010001","000000000000010000","000000000000001001","000000000000001100","111111111111110110","000000000000110000","000000000000101111","000000000000011101","111111111111101100","111111111111111100","111111111111111010","000000000000100011","111111111111100010","111111111111110000","000000000000100110","000000000000001100","111111111111110010","111111111111111100","111111111111001000","000000000000101001","000000000000001000","111111111111111100","000000000000010011","111111111111111111","000000000000000110","111111111111001011","111111111111110101","111111111111111110","111111111111111000","000000000000001010","111111111111010101","111111111111100110","111111111111100110","000000000000000000","111111111111110001","111111111111110001","111111111111110110","000000000000010111","000000000000001011","111111111111101110","111111111111110000","000000000000011011","111111111111110111","111111111111110110","000000000000001101","000000000000000111","111111111111111101","111111111111011111","000000000000011010","111111111111111111","000000000000010101","111111111111111001"),
("111111111111101101","000000000000000111","111111111111010111","111111111111111111","000000000000010011","000000000000000011","111111111111101000","111111111111110110","000000000000010111","111111111111011011","111111111111101010","000000000000000100","111111111111111110","111111111111001011","111111111111101001","111111111111101101","000000000000010001","111111111111111001","111111111111111000","000000000000011011","111111111111111001","000000000000010110","000000000000000100","111111111111100101","000000000000001011","000000000000001111","111111111111101101","000000000000000011","000000000000001011","000000000000010001","000000000000001000","111111111111111100","000000000000010100","000000000000001100","111111111111101100","111111111111110010","000000000000010101","000000000000010011","111111111111100010","000000000000011011","000000000000010000","111111111111111100","111111111111111110","111111111111000101","000000000000100001","111111111111100101","111111111111101011","000000000000100010","000000000000001011","000000000000000101","000000000000000111","000000000000011100","000000000000001000","111111111111111011","000000000000001011","111111111111110110","111111111111111001","000000000000011000","111111111111101101","000000000000000100","000000000000000000","000000000000000000","111111111111101010","111111111111101101","111111111111111001","000000000000000011","000000000000010111","111111111111100101","111111111111010100","000000000000000101","111111111111111111","000000000000001001","000000000000101001","111111111111011101","000000000000011100","111111111111110001","111111111111111001","000000000000010101","111111111111100010","000000000000011001","111111111111101111","000000000000101110","000000000000100101","000000000000001110","111111111111111110","111111111111101010","111111111111001110","000000000000010101","111111111111100100","111111111111101011","000000000000000011","000000000000011001","111111111111110111","111111111111111010","111111111111011100","000000000000010001","000000000000000000","000000000000001010","000000000000011000","000000000000001001","000000000000010001","111111111111111001","000000000000000010","000000000000010001","111111111111010101","000000000000010000","111111111111110100","111111111111011011","000000000000001011","000000000000001101","111111111111111100","111111111111100010","000000000000000100","000000000000001011","000000000000001110","000000000000000000","111111111111111100","000000000000000101","000000000000011010","000000000000001100","000000000000000001","111111111111111110","111111111111011011","111111111110101100","111111111111111010","111111111111101000","111111111111111111","000000000000000001"),
("111111111111101100","000000000000000111","111111111111001100","111111111111110100","000000000000001000","000000000000001000","000000000000000000","111111111111010111","000000000000010100","111111111111111101","111111111111110001","111111111111101110","000000000000010110","111111111111011011","000000000000001100","111111111111110111","000000000000000101","111111111111111100","111111111111111010","000000000000001111","000000000000000111","000000000000010000","000000000000000110","111111111111101100","000000000000010110","000000000000010000","111111111111001010","000000000000001001","111111111111111011","000000000000001010","000000000000100010","000000000000001010","111111111111110011","111111111111110100","111111111111011011","000000000000001100","111111111111111011","000000000000000001","111111111111110000","000000000000011001","000000000000000101","000000000000001101","111111111111011001","111111111111000111","000000000000100000","111111111111110011","111111111111000111","000000000000011011","000000000000011000","111111111111111011","000000000000010100","000000000000011000","000000000000001111","000000000000000000","000000000000011010","111111111111111011","111111111111110011","111111111111110110","000000000000010001","111111111111110110","000000000000000011","000000000000001111","111111111111110101","000000000000001000","111111111111101000","111111111111110110","111111111111111111","111111111111100110","111111111111000100","000000000000000001","111111111111101110","111111111111110111","000000000000100110","111111111111011100","000000000000100101","111111111111100011","000000000000010101","000000000000000110","111111111111101100","000000000000000101","111111111111101100","000000000000010000","000000000000001100","111111111111111100","000000000000000100","111111111111101101","111111111111011100","000000000000000111","111111111111110111","111111111111010110","000000000000000111","000000000000000000","111111111111100100","111111111111111011","111111111111001010","000000000000000111","111111111111110101","000000000000000011","000000000000011110","000000000000000100","000000000000001011","111111111111110011","000000000000000100","000000000000010010","000000000000000001","000000000000010011","111111111111011110","111111111111110101","111111111111011001","000000000000000000","111111111111111001","111111111111111110","111111111111111101","000000000000011000","000000000000000011","111111111111110100","000000000000000011","111111111111110101","111111111111101001","111111111111110111","111111111111111101","000000000000001110","111111111111100111","111111111110101011","111111111111011011","111111111111111000","000000000000000110","111111111111110000"),
("111111111111111101","000000000000010011","111111111111001101","000000000000010010","000000000000000000","000000000000000100","000000000000011110","111111111111001000","111111111111111111","111111111111100110","000000000000010001","111111111111111101","000000000000001110","111111111111101001","111111111111110011","000000000000000101","000000000000010110","000000000000010011","000000000000010011","000000000000011010","111111111111101101","000000000000010000","000000000000010001","000000000000000010","111111111111101100","000000000000010110","111111111111011100","111111111111111011","000000000000010100","111111111111110010","111111111111111011","111111111111110100","000000000000000110","111111111111101010","111111111111101011","111111111111101100","111111111111111010","000000000000000111","111111111111100100","111111111111110101","111111111111100101","111111111111111001","111111111111010110","111111111111001010","000000000000010000","000000000000000000","111111111111100101","111111111111100000","111111111111100100","111111111111110111","000000000000100100","000000000000000011","111111111111111100","111111111111011101","000000000000001101","000000000000000011","111111111111111101","000000000000000011","000000000000000100","111111111111111101","000000000000010000","000000000000011111","000000000000000100","000000000000000001","111111111111011000","111111111111111011","000000000000010010","000000000000001001","111111111110101101","000000000000000110","111111111111111101","000000000000010110","000000000000011010","111111111111100101","000000000000000001","111111111111011111","111111111111111111","000000000000001001","000000000000010100","111111111111111110","111111111111100110","111111111111111011","000000000000011010","000000000000001110","000000000000000111","111111111111011100","111111111110111010","000000000000001000","111111111111111001","111111111111100101","000000000000010010","000000000000000101","111111111111110101","000000000000000111","111111111111010100","111111111111011010","111111111111101110","111111111111110101","000000000000111011","000000000000000000","000000000000011000","111111111111010100","000000000000000101","111111111111101001","000000000000011001","000000000000010110","111111111111010101","111111111111101111","111111111111001001","000000000000010100","111111111111111000","000000000000000001","111111111111111100","111111111111111000","111111111111101011","000000000000011101","111111111111111010","111111111111110101","111111111111011100","000000000000001000","000000000000001001","111111111111110111","111111111111011010","111111111111001011","111111111111101010","111111111111110101","000000000000000100","111111111111110100"),
("111111111111111100","000000000000010011","111111111111011010","000000000000001111","111111111111101000","111111111111110110","000000000000101010","111111111111001110","000000000000001100","000000000000000000","000000000000010100","111111111111101001","000000000000010100","111111111111001110","111111111111101110","111111111111110010","111111111111111110","111111111111111110","000000000000010111","000000000000001000","000000000000000010","000000000000011000","000000000000011111","000000000000001100","000000000000001101","000000000000010000","111111111111111100","111111111111111101","111111111111111111","111111111111101010","000000000000010100","111111111111111100","000000000000000011","111111111111100111","000000000000010111","111111111111101110","000000000000000100","111111111111111110","111111111111010000","000000000000001001","111111111111101010","111111111111111100","111111111110101100","111111111111010111","000000000000010010","111111111111111001","000000000000000000","111111111111110111","000000000000000001","000000000000000000","000000000000110010","000000000000011101","000000000000011101","111111111111111010","000000000000011101","000000000000001000","000000000000001110","000000000000010110","000000000000000001","111111111111111101","000000000000011000","000000000000010010","000000000000100000","000000000000011001","111111111111000001","000000000000000000","000000000000000101","000000000000001111","111111111110111110","000000000000000001","111111111111101111","000000000000001110","000000000000010011","111111111111010110","111111111111110010","111111111111101010","000000000000000010","000000000000000100","000000000000000010","000000000000010110","000000000000001101","000000000000000000","000000000000001100","111111111111101000","111111111111111111","111111111111100110","111111111110110000","111111111111110111","111111111111101111","111111111111100010","000000000000000111","111111111111111010","111111111111110001","111111111111110111","111111111111010101","111111111111001101","111111111111101101","111111111111111001","000000000000101101","000000000000000101","000000000000001011","111111111111110110","000000000000010001","111111111111110011","000000000000011011","000000000000001001","111111111111011111","111111111111101001","111111111110110100","111111111111111101","111111111111111011","000000000000000101","000000000000000110","111111111111101100","000000000000000000","000000000000011011","111111111111101111","111111111111111111","111111111111010011","000000000000000000","000000000000011011","000000000000000001","111111111111011001","111111111111001111","000000000000001001","000000000000001000","111111111111110110","111111111111111000"),
("111111111111100111","000000000000110010","111111111110111100","000000000000010001","111111111111110011","111111111111110111","000000000000010011","111111111111100010","000000000000000010","000000000000000010","000000000000011100","111111111111111001","000000000000010001","111111111111111011","111111111111010010","111111111111111011","000000000000001111","000000000000000011","000000000000011000","000000000000000001","111111111111111101","000000000000000010","000000000000001110","000000000000010010","111111111111111000","111111111111111011","000000000000011001","000000000000000101","000000000000000000","111111111111100110","000000000000000100","000000000000001001","111111111111111001","111111111111111011","000000000000011101","000000000000000000","111111111111101100","000000000000000000","111111111111101001","000000000000001011","111111111111101111","000000000000001100","111111111111011100","000000000000010100","111111111111111101","111111111111101000","000000000000100011","000000000000000001","111111111111101011","000000000000001001","000000000000001001","111111111111110111","000000000000010111","111111111111100001","000000000000000110","111111111111110000","111111111111101111","111111111111111111","111111111111111010","000000000000001011","111111111111111001","000000000000011001","000000000000100010","000000000000001111","111111111111010100","000000000000000010","000000000000001010","000000000000000000","111111111111000011","111111111111110011","000000000000010100","000000000000011111","000000000000100101","111111111111010110","000000000000010101","111111111111100001","000000000000011000","000000000000000111","111111111111111100","111111111111111111","000000000000001011","111111111111100001","000000000000001000","111111111111110101","111111111111111101","111111111111100110","111111111110110010","000000000000001111","111111111111111101","000000000000001101","111111111111111110","111111111111111010","111111111111100110","000000000000100000","111111111111110101","111111111110110111","111111111111111111","111111111111111001","000000000000010010","000000000000010110","111111111111110010","111111111111100001","111111111111110111","000000000000000111","000000000000001001","000000000000000101","111111111111001111","111111111111110110","111111111110110100","000000000000000000","111111111111101110","000000000000000000","000000000000010111","111111111111110111","111111111111110000","000000000000001001","000000000000010111","111111111111101001","111111111111001010","111111111111110110","111111111111110100","000000000000100000","111111111111110111","111111111110100001","111111111111111001","000000000000000010","000000000000010110","111111111111100100"),
("111111111111111110","000000000000110000","111111111111000011","000000000000010001","111111111111111000","111111111111111110","000000000000001001","111111111111111101","000000000000000111","111111111111110111","000000000000100010","111111111111111011","000000000000011100","111111111111111101","111111111111000000","000000000000001011","000000000000010101","111111111111110010","000000000000100111","111111111111111010","000000000000000011","111111111111111101","000000000000100110","000000000000010110","000000000000000001","000000000000010010","000000000000010110","000000000000001010","111111111111011101","111111111111011001","000000000000001101","000000000000000001","000000000000011001","000000000000000000","000000000000010010","111111111111101001","111111111111100111","111111111111110100","111111111111101100","111111111111101111","111111111111010010","000000000000000000","000000000000011000","000000000000110000","000000000000001111","111111111111011000","000000000000100000","111111111111110010","111111111111110001","111111111111101110","111111111111101001","000000000000001101","000000000000001110","111111111111010000","000000000000011110","111111111111110100","111111111111110110","000000000000000100","111111111111111100","000000000000001110","000000000000001110","000000000000010010","111111111111111101","000000000000001001","111111111111100100","000000000000001100","000000000000010110","000000000000010101","111111111111001000","111111111111010111","000000000000001011","000000000000000000","000000000000100101","000000000000000000","111111111111111001","111111111111111110","000000000000011010","000000000000001101","111111111111011101","000000000000000101","000000000000000001","000000000000000110","000000000000001101","111111111111100100","111111111111110000","111111111111110101","111111111110110000","000000000000000111","000000000000000100","000000000000000001","111111111111100010","111111111111100011","000000000000000111","000000000000100100","000000000000001010","111111111111100100","111111111111111000","000000000000000111","000000000000011010","000000000000001101","000000000000001100","111111111111101111","000000000000000001","111111111111111010","000000000000100000","000000000000001111","111111111111100011","000000000000011011","111111111110110010","111111111111011110","111111111111111010","000000000000011001","000000000000011000","111111111111110001","111111111111100010","000000000000001101","000000000000011011","111111111111101001","111111111111001011","111111111111101011","000000000000001101","000000000000011011","000000000000000100","111111111110111010","000000000000001000","000000000000000001","000000000000010011","111111111111110111"),
("111111111111110110","000000000000100000","111111111111000010","111111111111110110","000000000000000000","000000000000000101","111111111111100000","000000000000001100","111111111111100010","000000000000000111","000000000000110001","111111111111100001","000000000000000011","000000000000000111","111111111110111111","111111111111111010","000000000000000111","111111111111100000","000000000000100000","111111111111111001","111111111111101110","000000000000000100","000000000000010011","000000000000000110","111111111111100000","000000000000001011","000000000000010100","000000000000010011","111111111111011001","111111111111101100","111111111111111100","111111111111101101","000000000000000011","111111111111110011","000000000000101111","111111111111010000","000000000000000000","111111111111110101","111111111111101001","111111111111110100","111111111111011000","000000000000010111","000000000000011000","000000000000011110","000000000000010111","111111111111011000","000000000000011110","111111111111101110","111111111111110101","111111111111110001","111111111111100100","111111111111110110","000000000000000001","111111111111011000","000000000000001100","111111111111101000","111111111111111011","000000000000000100","111111111111111011","111111111111110111","111111111111110111","000000000000011001","000000000000010111","111111111111110100","111111111111100010","111111111111110110","111111111111111101","111111111111111010","111111111111000010","111111111111011101","111111111111110110","111111111111111000","000000000000010001","111111111111010011","111111111111100000","111111111111111010","000000000000011100","000000000000000111","111111111111100111","111111111111110001","111111111111111001","000000000000001011","000000000000001010","111111111111110001","111111111111010110","111111111111100010","111111111111001110","000000000000010011","000000000000011010","111111111111101100","111111111111100001","111111111111010110","000000000000000010","000000000000001101","000000000000011100","111111111111000000","000000000000001100","111111111111111001","000000000000001101","000000000000000000","000000000000000011","000000000000001101","111111111111100010","111111111111011100","000000000000000101","000000000000010101","111111111111101000","000000000000101111","111111111111011111","111111111111011011","111111111111011101","000000000000001001","111111111111111000","000000000000000101","111111111111010101","000000000000011101","111111111111111001","111111111111100111","111111111111101001","111111111111101100","000000000000000011","000000000000010001","000000000001000000","111111111111011011","000000000000010000","000000000000010100","000000000000000001","111111111111110011"),
("000000000000000101","000000000000000000","111111111111011011","000000000000001001","111111111111110000","111111111111111001","000000000000000101","000000000000100100","111111111111010010","111111111111111111","000000000000101001","111111111111111011","000000000000010010","000000000000100100","111111111111101011","111111111111111010","000000000000000000","111111111111111111","000000000000000101","000000000000010010","111111111111111111","111111111111101011","000000000000001100","000000000000001010","111111111111111111","000000000000000011","000000000000001110","111111111111110101","111111111111110010","000000000000001100","111111111111111000","000000000000000010","000000000000001001","000000000000001010","000000000000001111","111111111111000110","000000000000000111","111111111111101011","111111111111011110","111111111111111000","111111111111011101","111111111111111100","000000000000110110","000000000000010100","111111111111110110","111111111111101000","000000000000100101","111111111111110101","000000000000001001","111111111111101001","111111111111100010","111111111111110111","111111111111111001","111111111111010000","000000000000010010","111111111111111100","111111111111111001","000000000000001000","111111111111111100","111111111111111110","000000000000000000","000000000000101110","000000000000000110","000000000000000000","111111111111110010","000000000000001011","000000000000001000","000000000000000000","111111111111010010","000000000000000001","000000000000000011","111111111111111100","000000000000111111","111111111111101001","111111111111100111","000000000000001000","000000000000010110","111111111111111100","111111111111111011","000000000000011000","111111111111110111","000000000000000110","111111111111110010","000000000000001001","111111111111111110","111111111111100001","111111111110100100","000000000000100001","000000000000001010","000000000000000000","111111111111100011","111111111111100110","000000000000010011","000000000000010100","000000000000010000","111111111111001010","000000000000001011","111111111111111000","000000000000101010","000000000000010100","111111111111101010","000000000000100010","111111111111100101","111111111111100110","000000000000000000","111111111111110001","111111111111100111","000000000000101100","111111111111000011","111111111111110001","111111111111100111","111111111111111111","000000000000001111","111111111111110001","111111111111010101","000000000000011000","000000000000010101","111111111111111111","111111111111100000","000000000000000000","000000000000001010","111111111111111111","000000000001001011","000000000000000000","111111111111111100","000000000000010011","111111111111110100","111111111111101110"),
("111111111111111001","111111111111110101","111111111111110011","000000000000000010","000000000000001010","000000000000011000","000000000000001101","000000000000010001","111111111111111111","111111111111111000","000000000000101011","111111111111110100","000000000000000001","000000000000011100","111111111111111010","000000000000010101","111111111111111100","111111111111100110","000000000000010000","000000000000010001","000000000000001000","111111111111001001","111111111111101111","111111111111111010","111111111111110100","000000000000001001","000000000000000000","111111111111110011","111111111111110101","000000000000011001","111111111111111001","000000000000010010","000000000000001011","000000000000000101","000000000000100011","111111111111001111","111111111111111111","000000000000010000","111111111111011111","000000000000001110","111111111111100110","111111111111111100","000000000000100001","000000000000011100","111111111111111100","000000000000011011","111111111111111110","000000000000011001","111111111111111111","111111111111100001","111111111111111111","111111111111110110","111111111111100001","111111111111110010","000000000000001110","111111111111111101","111111111111101111","111111111111111001","111111111111111100","000000000000000110","111111111111110101","000000000000101100","000000000000001001","111111111111111100","000000000000001101","111111111111101011","000000000000000000","000000000000001011","111111111111001001","000000000000001001","111111111111111010","111111111111111100","000000000000101001","000000000000001000","111111111111110000","000000000000000010","000000000000000101","000000000000001000","000000000000010010","000000000000010100","111111111111110000","111111111111111001","111111111111110100","000000000000001001","000000000000001011","000000000000000000","111111111110011111","000000000000000011","111111111111111111","111111111111111111","111111111111101011","111111111111011111","111111111111110111","000000000000000101","000000000000001001","111111111111100001","000000000000000101","111111111111111011","000000000000100010","000000000000001011","111111111111101100","000000000000111010","111111111111100111","111111111111110111","111111111111110110","000000000000010010","111111111111101111","000000000000011000","111111111111010010","111111111111110111","111111111111101001","000000000000001001","000000000000000001","000000000000000011","000000000000000011","000000000000010001","000000000000000011","000000000000011101","111111111111101101","000000000000000100","111111111111111111","111111111111110101","000000000000011000","000000000000100100","000000000000000101","111111111111111010","111111111111110111","000000000000000010"),
("111111111111110110","111111111111011010","000000000000000011","000000000000000101","111111111111110110","000000000000000100","111111111111111111","111111111111110110","111111111111100001","111111111111110010","000000000000100101","111111111111100000","000000000000000000","111111111111011111","000000000000110111","000000000000000000","000000000000010001","111111111111100101","111111111111110101","000000000000001111","000000000000000000","111111111110111011","111111111111100100","111111111111110001","000000000000010001","111111111111110011","111111111111011111","000000000000000111","000000000000010110","111111111111111111","000000000000001001","000000000000000111","111111111111100111","000000000000010010","111111111111110000","111111111111110111","000000000000010111","000000000000001010","000000000000010101","000000000000000011","000000000000001111","111111111111111100","000000000000001111","000000000000000101","111111111111111111","000000000000100101","000000000000011001","000000000000000100","111111111111111000","000000000000001111","111111111111110101","000000000000001000","111111111111011100","000000000000001011","000000000000010110","000000000000001101","111111111111111011","111111111111111110","000000000000001000","111111111111110100","000000000000000000","000000000000001101","111111111111111100","111111111111101100","000000000000010111","000000000000000000","000000000000100001","000000000000000001","111111111111011100","000000000000010000","000000000000000001","000000000000001010","000000000000010111","000000000000001011","000000000000010011","000000000000011101","000000000000010000","111111111111111011","000000000000000101","000000000000010110","000000000000000010","111111111111100111","000000000000100111","111111111111101110","000000000000000010","000000000000000000","111111111111011000","000000000000010010","000000000000001101","111111111111111100","000000000000100100","111111111111010101","000000000000000111","000000000000001001","111111111111101100","000000000000000110","111111111111101001","111111111111110100","000000000000001111","000000000000001011","000000000000001111","000000000000000110","111111111111111000","111111111111101101","111111111111011011","111111111111100011","000000000000000000","111111111111111110","111111111111100000","000000000000001110","000000000000000000","111111111111111010","111111111111110110","111111111111110011","111111111111101111","000000000000001010","000000000000010011","000000000000000100","111111111111111110","111111111111111111","111111111111111101","111111111111011101","000000000000001011","000000000000101001","000000000000011001","111111111111100100","111111111111110000","111111111111111000"),
("111111111111110010","111111111111010100","000000000000011000","111111111111110011","000000000000000101","000000000000100100","000000000000001011","000000000000001111","111111111111101001","111111111111011011","000000000000011111","111111111111101010","000000000000011010","111111111110111110","000000000000100101","111111111111110110","000000000000011011","000000000000001000","000000000000010100","000000000000001110","111111111111111101","111111111111000111","000000000000001011","111111111111101101","111111111111100111","111111111111111000","111111111111101010","111111111111111110","000000000000001100","000000000000001010","000000000000000100","000000000000001000","111111111111110010","000000000000000010","111111111111110110","000000000000000011","000000000000010111","000000000000001011","000000000000001101","000000000000000111","000000000000011110","111111111111101001","000000000000010010","111111111111111101","000000000000001101","000000000000001100","000000000000011110","111111111111111110","111111111111111000","111111111111110001","000000000000000000","111111111111101100","111111111111010001","000000000000000101","000000000000010111","000000000000001110","000000000000001010","111111111111111101","111111111111101110","000000000000000011","000000000000000110","000000000000000001","000000000000010000","111111111111110010","111111111111011011","111111111111110100","000000000000100011","000000000000011000","111111111111110001","111111111111110101","111111111111111010","000000000000000011","000000000000100111","111111111111101001","000000000000010110","000000000000100100","111111111111110011","111111111111110001","111111111111111101","000000000000010010","000000000000010111","111111111111100111","000000000000011000","111111111111010110","000000000000001110","000000000000011101","111111111111110111","000000000000001011","000000000000000101","000000000000000011","000000000000111010","111111111111101111","111111111111101100","111111111111101001","000000000000001001","111111111111111011","000000000000010001","111111111111100010","000000000000100111","111111111111111110","000000000000011101","111111111111111101","000000000000001110","000000000000001101","111111111111101100","111111111111110011","000000000000000101","000000000000000011","000000000000000111","000000000000001111","111111111111111111","111111111111111111","000000000000000000","000000000000010000","000000000000000110","000000000000010010","111111111111110101","000000000000001010","000000000000001010","000000000000000010","000000000000001010","000000000000001000","111111111111110111","000000000000111000","000000000000010001","111111111111100111","000000000000000000","000000000000000111"),
("000000000000000000","111111111111100100","000000000000010011","000000000000000110","000000000000001100","000000000000000000","111111111111111011","111111111111001001","000000000000000101","111111111111111001","000000000000000000","111111111111101110","000000000000011000","111111111111001011","000000000000001101","111111111111111110","000000000000010011","000000000000010100","000000000000000000","000000000000001100","111111111111111000","111111111111100101","000000000000011011","000000000000001000","111111111111111100","000000000000010111","111111111111111011","000000000000000010","000000000000011110","000000000000000101","111111111111110110","000000000000000110","000000000000010000","111111111111110101","111111111111110001","000000000000011110","111111111111110111","000000000000001101","000000000000010010","000000000000000001","000000000000101001","111111111111101000","000000000000000011","111111111111111100","000000000000010001","111111111111110011","000000000000000000","000000000000010100","000000000000000001","000000000000000111","111111111111110100","111111111111111111","111111111111011111","000000000000001111","111111111111101110","111111111111111011","000000000000001100","000000000000000000","111111111111111100","111111111111110100","000000000000010110","111111111111101010","000000000000010000","111111111111111000","111111111111001110","111111111111110101","000000000000100011","000000000000011001","111111111111110010","111111111111101101","111111111111111111","000000000000010010","111111111111110111","000000000000001011","000000000000001001","000000000000010100","111111111111111111","000000000000010000","111111111111111111","111111111111101001","000000000000001001","000000000000001111","000000000000101001","111111111111100011","000000000000001101","111111111111111001","000000000000100001","000000000000000101","000000000000000001","111111111111111111","000000000000011111","111111111111110001","000000000000000011","000000000000000000","111111111111101110","000000000000001000","000000000000001110","111111111111011010","000000000000101011","111111111111110010","000000000000010110","000000000000001100","000000000000100000","000000000000010001","111111111111110010","111111111111101110","111111111111110100","000000000000001000","000000000000000011","000000000000000110","111111111111101011","000000000000001110","000000000000000100","000000000000000000","111111111111111100","000000000000010000","000000000000010001","000000000000010000","000000000000000110","000000000000001001","111111111111111101","000000000000001001","111111111111010001","000000000000011110","000000000000001001","000000000000000001","000000000000000000","000000000000100001"),
("111111111111110110","111111111111111110","111111111111101110","111111111111111101","111111111111111000","000000000000000111","111111111111101000","111111111111010101","000000000000001000","000000000000100001","000000000000001101","000000000000000001","111111111111110010","111111111111101010","000000000000000101","000000000000010011","111111111111111010","000000000000011011","000000000000010000","000000000000010110","111111111111101011","000000000000100000","000000000000011010","111111111111110001","000000000000001001","000000000000001001","111111111111111001","111111111111110100","111111111111111101","000000000000000100","000000000000011001","000000000000010101","000000000000001011","000000000000000001","111111111111100001","111111111111111010","000000000000001001","000000000000001010","111111111111110011","000000000000010111","000000000000011010","000000000000000000","111111111111111011","000000000000000010","000000000000000000","111111111111110000","000000000000011011","000000000000100100","000000000000000001","000000000000001100","111111111111100000","000000000000001110","111111111111111011","000000000000001001","111111111111110000","111111111111110110","000000000000100100","000000000000000110","000000000000000010","111111111111111011","000000000000000100","000000000000001000","000000000000000100","111111111111111001","111111111111000100","111111111111111111","111111111111110101","000000000000010111","111111111111110101","111111111111101000","000000000000011010","000000000000001001","111111111111110111","111111111111111101","000000000000000100","111111111111110100","000000000000000000","000000000000000001","000000000000000001","111111111111101110","000000000000000000","111111111111111010","000000000000011101","111111111111110101","000000000000000110","111111111111101001","000000000000011010","111111111111111111","000000000000000011","000000000000001000","000000000000010100","000000000000001111","111111111111110111","000000000000000101","000000000000001011","000000000000011111","000000000000000011","111111111111101101","000000000000010001","111111111111101011","000000000000000011","111111111111111011","000000000000011100","000000000000100101","111111111111100100","000000000000000101","111111111111101110","000000000000001001","111111111111111010","111111111111111110","111111111111111111","000000000000101101","000000000000011010","000000000000011001","000000000000100011","111111111111111000","000000000000011100","111111111111111100","000000000000011100","000000000000000101","111111111111101000","111111111111110001","111111111111011111","000000000000100101","111111111111111101","111111111111101110","000000000000000101","111111111111111011"),
("111111111111111111","000000000000101001","111111111111110001","111111111111111011","111111111111110100","000000000000011001","111111111111110101","111111111111100110","111111111111101010","111111111111101010","000000000000000000","000000000000100000","000000000000000000","111111111111011001","111111111111111011","111111111111110111","111111111111110001","000000000000001110","111111111111111100","000000000000001000","000000000000001000","000000000000010011","000000000000010110","111111111111110001","111111111111110011","000000000000011111","000000000000010011","000000000000000110","111111111111100110","000000000000101001","000000000000000000","111111111111111101","000000000000010110","000000000000001010","000000000000000101","000000000000000111","111111111111101011","000000000000001101","000000000000010111","111111111111111010","111111111111110010","111111111111011010","000000000000010010","000000000000010110","000000000000100010","000000000000000101","000000000000011011","000000000000010000","111111111111111100","111111111111111100","111111111111101111","111111111111111110","111111111111110010","000000000000000011","000000000000000100","111111111111110101","000000000000100000","000000000000001111","000000000000001001","111111111111101101","000000000000100001","111111111111111101","000000000000100011","111111111111101000","111111111111001100","111111111111101010","111111111111101101","000000000000000101","000000000000000100","111111111111111010","111111111111111110","000000000000010000","000000000000000011","000000000000001000","000000000000010001","000000000000011010","111111111111110110","111111111111110010","111111111111101010","111111111111010110","000000000000001011","000000000000100010","000000000000001001","111111111111100111","000000000000100001","111111111111101110","111111111111111010","000000000000000110","111111111111111111","000000000000100000","000000000000001110","000000000000011000","111111111111101010","000000000000001111","111111111111110000","111111111111110110","111111111111110101","000000000000001010","000000000000000110","111111111111101111","000000000000010011","111111111111110010","000000000000100000","000000000000011010","111111111111110000","111111111111110001","111111111111101011","000000000000000011","111111111111101001","111111111111011001","111111111111111101","000000000000011110","111111111111111110","000000000000001010","000000000000000101","111111111111101101","000000000000010101","111111111111101011","000000000000000000","000000000000000010","111111111111111001","111111111111111011","111111111111111000","000000000000010100","000000000000010010","000000000000001001","000000000000001001","000000000000011011"),
("000000000000000000","000000000000101000","111111111111100101","000000000000000000","000000000000000110","000000000000001101","111111111111100001","000000000000011101","111111111111101111","111111111111111111","111111111111111011","000000000000010110","111111111111111011","111111111111110011","111111111111101110","000000000000000110","111111111111110000","000000000000011000","000000000000011001","111111111111111101","000000000000000110","000000000000001100","000000000000010110","000000000000000000","000000000000001011","000000000000000000","111111111111100111","111111111111111110","000000000000011010","111111111111110011","000000000000010011","000000000000000110","111111111111111110","000000000000000101","000000000000001101","000000000000000010","111111111111111000","000000000000000111","111111111111101101","000000000000000101","000000000000001110","111111111111110100","111111111111111000","000000000000010111","000000000000000100","111111111111111000","000000000000001000","000000000000011110","000000000000010001","000000000000001111","111111111111110001","000000000000001010","111111111111101011","000000000000100100","000000000000000011","000000000000000010","000000000000010001","000000000000000100","000000000000001101","111111111111101100","000000000000001101","111111111111111001","000000000000011001","111111111111101011","111111111111010111","000000000000001011","111111111111000001","000000000000010100","000000000000010110","000000000000000011","111111111111111111","000000000000011111","111111111111110110","111111111111111110","000000000000100101","000000000000010100","000000000000000100","111111111111111111","111111111111110000","111111111111100011","111111111111100010","000000000000001100","000000000000100001","111111111111100110","000000000000010011","111111111111100011","111111111111100011","000000000000000101","111111111111111001","111111111111111010","111111111111101010","000000000000000011","111111111111011111","000000000000001011","000000000000010101","111111111111011010","111111111111101000","111111111111110110","111111111111101100","000000000000010001","000000000000001110","111111111111111101","000000000000001110","000000000000011110","111111111111101100","111111111111101000","111111111111101100","111111111111100101","111111111111101110","111111111111111001","111111111111111110","111111111111111110","111111111111111100","111111111111110000","111111111111111000","111111111111110100","000000000000001000","111111111111111111","111111111111110011","000000000000001001","000000000000001010","000000000000000101","111111111111101110","000000000000001000","111111111111110011","000000000000010111","000000000000000000","000000000000001110"),
("000000000000001100","000000000001000000","000000000000000101","000000000000000000","111111111111110110","000000000000010001","111111111111111011","000000000000100110","111111111111101100","000000000000000000","000000000000001000","000000000000111011","111111111111100111","111111111111101110","111111111111010110","000000000000001111","000000000000000100","000000000000010000","111111111111111011","000000000000001110","000000000000000000","111111111111101001","000000000000001111","111111111111111000","000000000000001100","000000000000000000","111111111111110100","111111111111101010","000000000000010101","111111111111110100","000000000000000101","111111111111111001","111111111111100100","111111111111111110","000000000000000000","000000000000011000","000000000000001100","111111111111110111","000000000000000000","000000000000001010","111111111111111111","000000000000000001","111111111111110010","111111111111111100","000000000000010010","111111111111111011","000000000000000000","000000000000100101","000000000000011010","111111111111100111","111111111111101100","111111111111101101","000000000000000110","000000000000100011","000000000000001111","111111111111110010","111111111111100000","111111111111110111","000000000000001011","000000000000010001","000000000000000010","111111111111110100","111111111111111110","111111111111011111","111111111111100110","111111111111111110","111111111110110001","000000000000001110","000000000000011001","111111111111111111","111111111111101110","111111111111111011","111111111111010101","000000000000010100","000000000000000010","000000000000001101","000000000000000011","111111111111111111","111111111111100110","111111111111111111","111111111111011011","000000000000000000","000000000000010000","111111111111101100","000000000000010001","111111111111010101","000000000000000000","000000000000000110","000000000000000010","000000000000010010","111111111111111011","000000000000001011","111111111111110001","000000000000001101","000000000000010110","111111111111000101","111111111111101101","111111111111101111","111111111111100100","000000000000001000","000000000000001000","111111111111101100","111111111111011101","111111111111111100","111111111111100011","111111111111110010","111111111111110001","111111111111001100","111111111111110000","111111111111101010","111111111111111011","111111111111111000","000000000000000111","111111111111110011","111111111111100000","111111111111100011","111111111111100111","111111111111101101","111111111111001000","000000000000001001","000000000000001111","111111111111110011","000000000000000100","111111111111101101","111111111111101001","111111111111110111","000000000000001110","111111111111110111"),
("000000000000011001","000000000000100001","000000000000000000","111111111111110001","111111111111111101","000000000000000111","111111111111110001","000000000000000000","111111111111111010","000000000000000110","111111111111101110","000000000000011011","111111111111100011","111111111111111100","111111111111001100","000000000000000000","000000000000010101","000000000000000111","111111111111100001","000000000000000111","000000000000000110","111111111111110001","000000000000001111","111111111111101010","111111111111011000","000000000000001111","000000000000001000","111111111111011001","000000000000000001","111111111111001000","000000000000000101","111111111111110101","111111111111111100","000000000000000101","111111111111111110","000000000000001000","111111111111101110","000000000000000100","111111111111110001","000000000000010000","000000000000100110","111111111111111011","000000000000001000","111111111111101100","000000000000000100","111111111111110101","111111111111100010","111111111111111100","000000000000001110","111111111111111101","000000000000001001","111111111111110010","111111111111111011","000000000000010000","000000000000001110","111111111111110101","111111111111101010","111111111111100001","111111111111110001","111111111111111100","111111111111001101","000000000000000100","000000000000011001","111111111111110000","111111111111111100","111111111111101111","111111111110011111","111111111111110010","000000000000100111","111111111111100011","000000000000001010","111111111111110001","111111111110101011","000000000000000000","000000000000000000","000000000000000010","000000000000010011","111111111111011001","111111111111111011","000000000000000110","111111111111011010","111111111111111001","000000000000000010","111111111111010100","000000000000011001","111111111111100010","111111111111101111","000000000000000010","111111111111111001","000000000000011100","000000000000000110","000000000000001010","000000000000000100","000000000000001100","111111111111110111","111111111111000001","111111111111111010","111111111111110001","111111111111010111","111111111111110100","000000000000010011","111111111111101110","111111111111010011","000000000000011101","111111111111011010","000000000000001101","111111111111110101","111111111111100000","000000000000000000","111111111111111010","000000000000000001","000000000000001001","000000000000011010","000000000000001001","111111111111100111","111111111111100010","111111111111110111","111111111111110101","111111111111100011","000000000000010101","000000000000001110","111111111111111001","111111111111111010","111111111111011001","000000000000001100","111111111111111000","000000000000001001","000000000000001001"),
("000000000000100101","000000000000010000","111111111111011111","000000000000010011","111111111111010100","000000000000011001","000000000000011000","000000000000001011","000000000000010010","111111111111101111","111111111111101000","000000000000100010","000000000000000000","111111111111111001","111111111111100101","000000000000000110","000000000000000000","000000000000000101","111111111111011100","111111111111110101","000000000000010011","111111111111110011","000000000000100001","111111111111110011","111111111111111110","000000000000000000","111111111111110101","111111111111101001","000000000000000001","111111111111011110","000000000000001011","111111111111110110","111111111111101100","000000000000001111","000000000000000000","111111111111110100","000000000000000111","000000000000011000","111111111111110001","111111111111110100","000000000000010100","111111111111101000","000000000000010110","000000000000000101","111111111111101100","111111111111110010","111111111111111001","000000000000011010","111111111111100001","111111111111110011","000000000000101000","000000000000001111","000000000000001101","000000000000000000","000000000000011001","111111111111101101","111111111111100001","111111111111110110","111111111111111101","000000000000001010","111111111111010001","111111111111111011","000000000000000000","000000000000000111","000000000000001101","111111111111011010","111111111110111010","111111111111111010","000000000000001010","111111111111111010","000000000000101100","111111111111111011","111111111111011110","000000000000000111","000000000000000000","111111111111111111","000000000000000000","111111111111011010","111111111111010100","111111111111111111","111111111111101111","000000000000001000","000000000000010101","111111111110111010","000000000000101101","111111111111011010","111111111111110110","000000000000010101","000000000000000001","111111111111111010","111111111111111011","000000000000000100","111111111111101110","000000000000011010","111111111111111001","111111111111100011","111111111111110110","111111111111101110","111111111111100000","111111111111101110","000000000000100100","000000000000001001","111111111111010101","000000000000010110","111111111111101101","000000000000100100","111111111111011001","111111111111110100","111111111111111100","111111111111101011","111111111111111100","111111111111111001","000000000000011010","000000000000001101","111111111111110110","000000000000011100","000000000000000100","000000000000011101","111111111111011110","000000000000001111","111111111111110001","000000000000010001","111111111111111111","111111111111010100","111111111111111011","000000000000001110","111111111111110111","111111111111111010"),
("000000000000101000","000000000000001111","111111111111100100","000000000000000001","111111111111100110","000000000000001101","000000000000000101","000000000000000101","000000000000011100","000000000000000000","111111111111101101","000000000000000111","000000000000010100","000000000000010010","111111111111100100","111111111111111101","000000000000001011","000000000000001110","111111111111011110","111111111111111101","000000000000010010","111111111111011010","111111111111101010","111111111111100001","111111111111110100","000000000000101111","000000000000001011","111111111111110110","111111111111101100","111111111111110100","000000000000010100","111111111111100110","111111111111110110","111111111111111101","111111111111110111","000000000000000011","111111111111101101","000000000000100001","111111111111011111","111111111111110001","000000000000010110","111111111111100100","000000000000001000","000000000000010100","111111111111111111","111111111111100100","000000000000000011","000000000000101011","111111111111011011","111111111111110100","000000000000101101","111111111111111110","111111111111111011","000000000000001110","000000000000011110","000000000000010110","111111111111011001","111111111111111000","111111111111010111","111111111111110100","111111111111001001","111111111111110011","000000000000100101","111111111111101010","111111111111111110","111111111111011111","111111111111100000","111111111111110111","111111111111111110","111111111111111001","000000000000100001","111111111111111001","111111111111100111","111111111111101110","000000000000001001","000000000000011111","000000000000000011","111111111111100010","111111111111100011","000000000000001000","111111111111101100","111111111111110011","000000000000100110","111111111110110011","000000000000100010","111111111110111110","111111111111101000","000000000000010100","000000000000010001","111111111111011101","000000000000000000","111111111111110101","111111111111111111","000000000000000000","111111111111101110","000000000000000011","000000000000001000","111111111111110100","111111111111011101","111111111111010011","000000000000011111","000000000000001000","111111111111011111","000000000000011001","111111111111110010","000000000000100011","111111111111010110","111111111111111000","111111111111011001","111111111111101000","000000000000000000","111111111111101001","000000000000010100","111111111111110101","111111111111101100","000000000000000010","000000000000000011","000000000000000001","111111111111011100","111111111111111101","111111111111101101","000000000000010110","000000000000010110","111111111111100110","000000000000001110","000000000000000100","111111111111111000","111111111111001000"),
("000000000000101111","000000000000011000","111111111111111101","000000000000001110","111111111111101001","000000000000001101","111111111111111000","111111111111110011","111111111111111100","111111111111110010","111111111111101011","000000000000010001","000000000000010010","000000000000010100","111111111111100101","111111111111110111","111111111111110110","000000000000100011","111111111111100100","111111111111111000","000000000000111011","111111111111110010","111111111111111100","111111111111110010","000000000000000010","000000000000001010","000000000000101100","111111111111101101","000000000000001000","111111111111010111","000000000000000100","111111111111110101","111111111111011101","111111111111111110","000000000000010101","111111111111111111","000000000000000000","000000000000000101","111111111111010000","111111111111101101","000000000000000001","111111111111110011","111111111111110001","000000000000000111","111111111111101010","111111111111100110","111111111111011110","000000000000110101","000000000000000101","111111111111011110","111111111111111011","000000000000000010","111111111111111111","000000000000100011","000000000000011001","000000000000001110","111111111111111011","000000000000010000","111111111111011111","000000000000001100","111111111111111001","000000000000001111","000000000000011011","000000000000001001","000000000000011110","111111111111100010","111111111111111100","111111111111011011","111111111111101110","111111111111100101","111111111111110110","000000000000011111","111111111111111110","111111111111111111","000000000000000000","111111111111110011","111111111111110011","111111111111100011","111111111111101000","111111111111100001","000000000000000000","111111111111110111","000000000000000111","111111111111010011","000000000000011011","111111111111000100","000000000000001010","000000000000001010","111111111111111110","111111111111100010","000000000000100100","000000000000000010","000000000000000101","111111111111111100","111111111111111011","111111111111101101","000000000000000000","111111111111100010","111111111111111010","111111111111101110","111111111111111111","000000000000010101","111111111111001101","000000000000011000","111111111111111001","000000000000001111","111111111111101111","111111111111110101","111111111111001111","111111111111011100","000000000000000110","111111111111101110","111111111111011101","111111111111101101","111111111111101000","111111111111110100","111111111111000101","000000000000010010","111111111111100111","000000000000000010","000000000000000000","000000000000100111","000000000000011011","111111111111101010","000000000000000001","000000000000000101","111111111111110001","111111111111011111"),
("000000000000100011","111111111111101000","000000000000001001","000000000000100000","000000000000010100","000000000000100000","000000000000000101","000000000000100000","000000000000011110","111111111111100100","000000000000101011","111111111111101000","000000000000100100","000000000000100101","111111111111100000","000000000000010000","000000000000000001","000000000000001011","111111111111000111","111111111111111010","000000000000011001","111111111111011000","111111111111100001","000000000000011010","111111111111111010","000000000000010101","000000000000000100","000000000000001011","000000000000011100","111111111111111101","000000000000101110","111111111111110110","111111111111101100","111111111111110000","000000000000100100","000000000000000110","000000000000000100","000000000000011110","111111111111111000","111111111111010110","111111111111100110","000000000000000100","000000000000100110","000000000000100001","111111111111000011","111111111111111101","111111111111100101","000000000000101011","111111111111000110","111111111111011001","111111111111101000","111111111111110100","111111111111110110","000000000000111001","000000000000011010","111111111111110000","000000000000000001","111111111111101010","111111111111000100","000000000000000000","000000000000000110","000000000000010100","000000000000011010","111111111111101011","000000000000000100","111111111111001011","000000000000011010","111111111111101001","111111111111110111","111111111111100011","000000000000011101","000000000000001100","000000000000100001","111111111111100001","000000000000001001","000000000000000110","000000000000000010","111111111111111001","111111111111010100","111111111111101111","000000000000000011","111111111111100001","000000000000001100","111111111111100011","000000000000100000","111111111111111100","000000000000011111","000000000000101010","111111111111100011","111111111111101101","111111111111111111","111111111111101011","111111111111111011","000000000001000100","111111111111001100","111111111111101101","111111111111110000","111111111111110010","000000000000001010","111111111111110010","000000000000001000","111111111111101111","111111111111010110","111111111111111001","000000000000000110","000000000000000000","111111111111100001","111111111111110100","111111111111011110","111111111111101110","111111111111111100","000000000000001010","111111111111100111","111111111111010010","111111111111000110","000000000000000000","111111111111011111","000000000000101001","000000000000000111","111111111111101001","000000000000011101","000000000000111110","000000000000000100","111111111111100101","000000000000100001","111111111111110100","111111111111111000","000000000000000011"),
("111111111111111111","111111111111001001","000000000000000010","000000000000000000","111111111111111110","000000000000110011","111111111111111000","000000000000100010","000000000000101011","111111111111000101","000000000000100010","111111111111011101","000000000000100010","000000000000000011","111111111111101001","000000000000100001","000000000000111000","000000000000101000","111111111111011010","000000000000001111","000000000000000010","111111111111101110","111111111111110001","000000000000000000","111111111111111001","000000000000101010","111111111111100101","000000000000001001","000000000000001101","111111111111101111","000000000000100100","111111111111100011","111111111111111100","111111111111011100","000000000000010101","111111111111111101","000000000000011011","000000000000100110","111111111111111100","111111111111011000","111111111111010000","111111111111110100","000000000000101000","000000000000110100","111111111111110000","000000000000001011","000000000000000111","111111111111111101","111111111111010111","111111111111111101","111111111111011101","000000000000000011","111111111111111110","000000000000000000","000000000000100101","000000000000011011","111111111111110100","111111111111111100","111111111111101100","111111111111101100","111111111111111010","000000000000101000","000000000000100110","000000000000100000","000000000000100000","111111111111011011","000000000000000010","111111111111100111","000000000000011110","111111111111011111","000000000000010111","000000000000000010","111111111111111111","000000000000010111","111111111111111000","000000000000011111","000000000000010110","111111111111111110","000000000000001100","111111111111111010","111111111111101101","000000000000001000","000000000000011111","000000000000010001","000000000000010110","111111111111101100","000000000000001110","000000000000001010","111111111111111011","000000000000000100","111111111111001111","111111111111110010","000000000000000111","000000000000001011","111111111111111110","000000000000000111","111111111111010011","111111111111111100","111111111111111011","111111111111011111","000000000000011100","111111111111111010","111111111111010111","000000000000000001","111111111111110101","000000000000000100","111111111111110000","111111111111111100","111111111111111101","111111111111100101","111111111111110111","000000000000011110","111111111111110101","111111111111111001","000000000000001011","000000000000000110","111111111111111011","000000000000001111","000000000000000000","000000000000010001","000000000000100111","000000000000110111","000000000000010111","000000000000100000","000000000000100001","111111111111101111","000000000000011010","000000000000000001"),
("000000000000000101","111111111111110111","111111111111110110","000000000000011000","000000000000011101","000000000000001100","000000000000001010","000000000000101011","111111111111111100","111111111111101010","000000000000010110","111111111111100001","000000000000011001","000000000000001100","111111111111100111","000000000000011101","000000000000001100","000000000000010000","000000000000000010","000000000000100010","000000000000011000","111111111111110110","000000000000010011","000000000000000101","111111111111110101","000000000000001001","111111111111110110","000000000000011010","000000000000011011","111111111111111100","000000000000000011","000000000000010010","111111111111111101","111111111111110010","000000000000011111","111111111111110110","000000000000001010","111111111111111000","111111111111111011","111111111111101010","111111111111010111","000000000000010011","000000000000011000","000000000000000001","111111111111111001","111111111111100011","000000000000000100","111111111111111111","111111111111101011","000000000000000000","111111111111110010","000000000000011011","111111111111110101","111111111111101000","000000000000010101","000000000000000100","111111111111101011","111111111111111011","000000000000001010","111111111111110000","000000000000000010","000000000000101010","000000000000001100","000000000000000100","000000000000010100","111111111111111001","111111111111101000","000000000000000000","111111111111110000","111111111111111011","111111111111101010","111111111111101110","000000000000100101","000000000000011101","111111111111100001","000000000000000110","000000000000000001","111111111111110011","000000000000000100","000000000000000001","111111111111100010","000000000000000000","111111111111101101","000000000000011110","000000000000000101","000000000000001011","111111111111110000","111111111111111010","000000000000000101","111111111111101001","111111111111101010","000000000000001001","000000000000000100","000000000000001101","111111111111110000","111111111111100101","111111111111101100","111111111111110100","111111111111011100","000000000000001100","000000000000101010","000000000000000000","111111111111101111","111111111111100010","000000000000000000","000000000000000101","111111111111100001","111111111111100101","000000000000010100","111111111111110011","111111111111011101","000000000000001010","111111111111110011","000000000000000011","111111111111101100","000000000000001110","000000000000000001","000000000000101100","000000000000001010","000000000000010010","000000000000000101","000000000000000011","000000000000011000","111111111111101111","000000000000010001","111111111111111100","000000000000011011","000000000000011001"),
("111111111111101110","111111111111110100","111111111111101101","000000000000001001","000000000000001111","000000000000000110","111111111111111101","111111111111111101","111111111111111110","111111111111110011","000000000000000010","000000000000001000","000000000000000011","111111111111111111","000000000000000100","111111111111110010","111111111111111000","000000000000000101","000000000000001101","000000000000010000","000000000000000011","000000000000001110","111111111111110100","111111111111111100","000000000000001100","111111111111111111","111111111111110000","111111111111111100","111111111111111011","111111111111110010","000000000000000111","000000000000010010","000000000000001101","111111111111110101","111111111111111111","000000000000000100","111111111111111011","111111111111111111","000000000000001011","000000000000001010","111111111111111101","000000000000000000","000000000000001111","111111111111111000","111111111111101111","111111111111110000","000000000000010011","111111111111101101","111111111111110010","111111111111111101","111111111111110010","111111111111111000","000000000000001000","000000000000000011","000000000000000010","000000000000000010","000000000000001011","111111111111110110","000000000000001110","000000000000001010","000000000000010011","000000000000000110","000000000000000111","000000000000000111","000000000000001000","000000000000001011","000000000000001100","000000000000001001","000000000000001100","111111111111110110","111111111111111001","111111111111111000","111111111111111000","111111111111111011","111111111111110001","000000000000000100","111111111111111010","111111111111111010","111111111111101110","000000000000000111","000000000000001101","111111111111111111","111111111111110100","111111111111111010","111111111111110001","111111111111111101","111111111111101100","111111111111110101","000000000000010001","000000000000010010","000000000000001101","111111111111101101","111111111111111111","000000000000001011","111111111111110100","000000000000010001","000000000000001100","000000000000001111","111111111111110101","000000000000010000","000000000000000011","111111111111111011","000000000000000010","111111111111101101","000000000000000000","111111111111111001","000000000000001000","111111111111110110","000000000000000111","000000000000010100","111111111111101110","000000000000010010","000000000000010001","111111111111110001","000000000000000001","111111111111101101","111111111111111000","000000000000001101","111111111111111010","000000000000001011","000000000000010000","111111111111110110","111111111111111111","111111111111110001","111111111111111011","000000000000001001","111111111111111101","000000000000001011"),
("000000000000000000","111111111111101011","000000000000000011","111111111111111010","000000000000000001","111111111111111011","111111111111111110","000000000000001111","111111111111110011","111111111111110100","000000000000000100","000000000000000100","000000000000001110","111111111111111111","000000000000000011","000000000000000100","111111111111111010","000000000000010011","111111111111111100","000000000000010101","111111111111110111","000000000000001000","111111111111111001","000000000000011011","000000000000000101","111111111111101000","000000000000001001","000000000000011101","111111111111111001","000000000000011001","111111111111110010","111111111111111001","000000000000011101","111111111111101100","000000000000000111","111111111111101111","111111111111110011","111111111111110110","111111111111110000","000000000000001110","111111111111110101","111111111111101010","000000000000010101","000000000000000101","000000000000000000","111111111111110011","111111111111111101","111111111111101000","000000000000011001","111111111111110000","000000000000011110","000000000000010000","111111111111111110","000000000000001000","000000000000001101","000000000000000010","000000000000000010","000000000000000000","000000000000010001","111111111111111000","111111111111111011","000000000000001010","111111111111111101","000000000000010101","000000000000000001","000000000000001111","000000000000011010","000000000000010010","000000000000001011","111111111111101110","111111111111111000","111111111111111101","000000000000000000","000000000000011100","000000000000001100","111111111111111111","111111111111110000","000000000000001101","111111111111101001","000000000000010110","111111111111110111","000000000000001110","111111111111101110","000000000000011010","000000000000010101","000000000000010000","111111111111100101","111111111111111100","000000000000001001","111111111111111011","000000000000001110","000000000000011011","111111111111110100","000000000000011000","000000000000010111","111111111111111101","000000000000011000","111111111111111001","111111111111110111","000000000000010001","111111111111111010","000000000000000000","000000000000001000","000000000000010100","111111111111110101","000000000000010010","111111111111101111","000000000000000001","000000000000000111","111111111111110101","000000000000001001","111111111111111110","111111111111110111","000000000000000011","000000000000001100","000000000000011010","000000000000000001","111111111111111100","000000000000001101","000000000000010101","111111111111100011","111111111111110100","000000000000001111","111111111111111101","000000000000001000","000000000000000010","000000000000001101","111111111111110111"),
("111111111111111000","111111111111110110","111111111111111101","111111111111110110","000000000000001000","000000000000001100","000000000000001001","000000000000000010","000000000000000100","111111111111110000","000000000000010110","000000000000011010","000000000000010011","111111111111100101","111111111111101000","000000000000011010","000000000000001001","000000000000000111","000000000000010011","000000000000010011","111111111111101111","111111111111111111","111111111111111001","111111111111010110","000000000000000000","000000000000011111","111111111111100110","111111111111110111","000000000000000110","111111111111111000","000000000000101101","111111111111110101","000000000000000000","000000000000000100","000000000000000100","111111111111110101","000000000000001001","000000000000100011","111111111111110110","111111111111111011","111111111111110100","000000000000011000","111111111111110001","111111111111101100","000000000000010001","111111111111111011","000000000000001111","000000000000001100","111111111111111011","111111111111101101","111111111111101011","000000000000011110","000000000000010110","000000000000000010","111111111111111010","000000000000010001","111111111111111010","111111111111100000","111111111111011001","111111111111110100","111111111111110110","000000000000010000","000000000000000000","000000000000001101","111111111111010100","111111111111111001","111111111111011001","000000000000000100","111111111111110100","111111111111111001","000000000000000111","111111111111100100","111111111111101001","111111111111011110","111111111111011110","000000000000001001","000000000000011001","111111111111111100","000000000000010110","000000000000010000","111111111111110000","000000000000001001","000000000000100011","111111111111111010","111111111111100111","000000000000000010","000000000000001111","111111111111101100","000000000000000110","111111111111100100","000000000000000001","111111111111100010","111111111111101000","111111111111101100","111111111111101101","000000000000000010","111111111111111011","000000000000011000","000000000000000011","111111111111101101","000000000000001001","111111111111111101","111111111111011100","000000000000001000","000000000000010110","000000000000001101","111111111111100111","111111111111101101","111111111111111111","111111111111110110","000000000000000101","000000000000101100","111111111111101011","111111111111111011","000000000000001000","111111111111110000","111111111111110010","000000000000100001","000000000000000001","111111111111100100","000000000000011100","000000000000010001","111111111111100110","111111111111110111","000000000000010000","000000000000010011","000000000000010101","111111111111111001"),
("000000000000000010","111111111111101000","111111111111110011","000000000000001010","000000000000001011","000000000000001100","111111111111100111","000000000000000011","000000000000010110","111111111111101010","000000000000011001","000000000000001010","000000000000101100","111111111111000001","111111111111100010","000000000000010000","000000000000101101","111111111111101000","000000000000100001","000000000000100001","111111111111011010","111111111111101101","111111111111111111","111111111111010111","111111111111010010","000000000000100111","111111111111110010","000000000000001111","000000000000110000","111111111111101111","000000000000000000","111111111111111000","000000000000010110","111111111111111100","000000000000000011","000000000000010001","111111111111110010","000000000000001010","111111111111111101","000000000000010101","000000000000000101","111111111111111101","111111111111101100","111111111111011010","000000000000100110","111111111111111011","000000000000001001","111111111111100110","111111111111101111","111111111111111011","000000000000010000","000000000001001000","111111111111011101","000000000000011000","000000000000011100","000000000000000000","111111111111011011","000000000000001000","111111111111011000","000000000000000000","111111111111110001","000000000000011001","000000000000100000","111111111111101101","111111111111111000","111111111111011000","111111111110111001","111111111111110001","111111111111110010","111111111111111101","111111111111111110","000000000000000100","111111111111000110","111111111111100100","000000000000100101","000000000000110000","000000000000001000","000000000000110001","000000000000000000","000000000000100110","111111111111101001","000000000000101000","000000000000101011","000000000000001111","111111111111111110","111111111111110111","000000000000000100","000000000000100111","111111111111110011","111111111111101001","111111111111100011","111111111111111011","111111111111101101","111111111111110001","111111111111010100","000000000000100000","111111111111101000","000000000000010000","000000000000010001","111111111111110100","111111111111111001","111111111111110010","111111111111111011","000000000000000101","111111111111101010","000000000000000110","111111111111011001","111111111111100011","000000000000101011","000000000000000011","111111111111100001","000000000000100111","000000000000010101","111111111111110111","000000000000000111","111111111111111111","111111111111111000","000000000000100101","111111111111101011","000000000000011011","000000000000100111","111111111111101011","111111111111111110","111111111110111100","000000000000111010","000000000000001110","000000000000100000","111111111111110011"),
("111111111111110100","111111111111101101","111111111111010111","000000000000001001","000000000000000110","000000000000000000","111111111111101111","000000000000001011","000000000000000111","111111111111011100","000000000000010010","111111111111110101","000000000000001110","111111111111010010","111111111111101110","000000000000010001","000000000000010001","111111111111110110","111111111111101101","000000000000000000","111111111111110010","000000000000010000","000000000000001000","111111111111010010","111111111111111101","000000000000010001","111111111111010010","000000000000001000","000000000000001000","000000000000000001","000000000000001000","000000000000010111","000000000000001111","000000000000011100","111111111111110101","000000000000100010","111111111111110001","000000000000011001","000000000000000000","000000000000000110","000000000000001000","111111111111110101","111111111111110001","111111111111101111","000000000000011110","111111111111101011","111111111111111010","000000000000000110","000000000000001100","111111111111110100","000000000000001101","000000000000100101","111111111111110110","000000000000010010","000000000000100010","111111111111100011","111111111111101100","000000000000000011","000000000000000111","111111111111111011","000000000000000001","000000000000001001","000000000000001011","000000000000000100","111111111111101110","111111111111110100","111111111111001111","000000000000000011","111111111111111000","000000000000001101","000000000000010010","000000000000011010","111111111111100001","111111111111101110","000000000000000000","111111111111111000","111111111111111001","000000000000011001","111111111111111000","000000000000010011","111111111111011011","000000000000111001","000000000000010101","000000000000011011","000000000000001111","000000000000000011","111111111111110010","111111111111110100","111111111111010101","111111111111010000","000000000000000100","000000000000011011","111111111111100100","111111111111110110","111111111111001001","000000000000110010","111111111111101100","111111111111111110","000000000000010110","111111111111100000","000000000000001110","111111111111011100","111111111111111000","000000000000010000","111111111111011011","000000000000000000","111111111111101111","111111111111100111","000000000000011101","000000000000010001","111111111111100110","000000000000100101","111111111111110111","000000000000001010","000000000000001011","000000000000000100","111111111111111101","000000000000001100","000000000000001010","000000000000011011","000000000000010101","111111111111111100","000000000000001010","111111111110111011","000000000000011101","000000000000001111","111111111111110010","000000000000000110"),
("111111111111101000","111111111111101100","111111111111010111","000000000000010110","111111111111101101","111111111111111011","000000000000010000","111111111111101100","000000000000010100","111111111111100100","111111111111110001","111111111111111110","000000000000001001","111111111111100010","111111111111111011","000000000000000010","000000000000000000","000000000000001101","111111111111101000","000000000000001111","111111111111110111","000000000000010101","111111111111111100","111111111111100110","000000000000011100","000000000000010101","111111111111000010","000000000000011010","111111111111010100","111111111111111111","000000000000011111","000000000000000101","000000000000110010","000000000000000011","111111111111110111","111111111111111001","000000000000001000","000000000000001101","111111111111111001","111111111111111101","000000000000000011","111111111111110110","111111111111110100","111111111110111111","000000000000010001","111111111111010110","111111111111011100","000000000000001001","111111111111110111","000000000000001100","111111111111111110","000000000000010000","000000000000001111","000000000000100100","000000000000011011","000000000000000111","000000000000010010","000000000000001001","000000000000001001","000000000000000011","000000000000001010","111111111111101111","111111111111101011","000000000000000101","111111111111101111","000000000000000100","000000000000000011","111111111111101110","111111111111001110","000000000000000100","111111111111110101","111111111111110110","000000000000000101","111111111111110000","000000000000010100","111111111111110000","000000000000001001","000000000000100001","111111111111100000","000000000000001011","000000000000000001","000000000000111101","000000000000001011","000000000000000000","111111111111111101","111111111111101001","111111111111111100","000000000000000010","111111111111100100","111111111111110010","111111111111111011","000000000000011101","111111111111100110","111111111111111000","111111111111100011","000000000000101111","000000000000000001","000000000000010001","000000000000001101","111111111111111000","111111111111110011","111111111111011110","000000000000000000","000000000000001010","111111111111111011","000000000000000101","111111111111110011","111111111111101110","000000000000010101","000000000000001110","000000000000000011","000000000000100100","000000000000000000","111111111111110011","000000000000000001","000000000000000001","000000000000000111","000000000000011011","000000000000010011","000000000000011100","000000000000000110","000000000000000100","111111111111011100","111111111110111010","111111111111100111","000000000000000101","000000000000011000","000000000000010000"),
("111111111111101001","111111111111111101","111111111110111010","000000000000010100","000000000000001000","000000000000001111","111111111111100100","111111111111101011","000000000000001100","111111111111101011","000000000000000100","111111111111101110","000000000000010110","111111111111100000","000000000000000011","111111111111111010","111111111111101100","000000000000101010","111111111111111111","000000000000001111","111111111111111110","000000000000000010","111111111111111101","000000000000000010","000000000000000010","000000000000000000","111111111111010101","111111111111110110","111111111111111001","111111111111111011","000000000000100100","000000000000100011","111111111111111010","000000000000000011","000000000000000111","000000000000000011","111111111111101001","000000000000000100","111111111111100000","000000000000010111","000000000000001001","111111111111101101","111111111111110101","111111111111010000","111111111111111111","000000000000010101","111111111111101110","111111111111110110","111111111111111001","000000000000010100","000000000000100000","000000000000011111","000000000000001100","000000000000001001","000000000000011000","000000000000001101","000000000000001101","111111111111110000","111111111111110010","111111111111101101","000000000000011001","000000000000000100","111111111111111011","111111111111101011","111111111110111011","000000000000000100","000000000000101011","111111111111100110","111111111111001100","111111111111101011","000000000000010010","000000000000100110","000000000000011110","111111111111101101","000000000000011110","111111111111111111","000000000000010001","000000000000010011","111111111111110110","111111111111101110","111111111111101011","000000000000011000","000000000000000000","111111111111111011","000000000000011101","111111111111100110","111111111111110110","000000000000011111","111111111111101111","111111111111111110","000000000000000101","111111111111111100","111111111111110011","111111111111100101","111111111111001011","000000000000010011","111111111111110011","111111111111101000","000000000000101011","000000000000001011","111111111111101010","111111111111100101","000000000000011101","000000000000001111","111111111111111111","000000000000010100","111111111111100001","111111111111101010","111111111111111010","111111111111101010","111111111111100100","000000000000000111","111111111111110010","000000000000010100","111111111111111001","000000000000000011","000000000000000110","000000000000000100","111111111111111100","000000000000001111","111111111111111100","000000000000001010","111111111111011010","111111111111001010","111111111111100111","111111111111111100","000000000000000100","111111111111111001"),
("111111111111101011","111111111111110011","111111111110111011","000000000000010100","000000000000000111","000000000000000001","000000000000000111","111111111111001111","000000000000011111","111111111111110101","000000000000100111","111111111111110011","000000000000011100","111111111111001000","111111111111110001","000000000000001101","000000000000001100","000000000000001101","000000000000001110","000000000000001110","111111111111110110","000000000000101001","000000000000001100","111111111111110000","111111111111101010","000000000000011111","000000000000001001","000000000000010110","000000000000011011","111111111111111011","000000000000001000","000000000000010001","111111111111101111","111111111111111110","000000000000000011","000000000000001001","111111111111111100","111111111111110110","000000000000000000","000000000000001000","000000000000000011","000000000000001010","111111111111001100","111111111111010000","000000000000010001","000000000000001000","111111111111110111","111111111111110100","111111111111111101","000000000000001010","000000000000100100","000000000000010111","111111111111110101","111111111111111110","000000000000000010","000000000000000000","111111111111100110","000000000000001111","111111111111101010","111111111111110010","000000000000010100","000000000000001101","000000000000011011","000000000000010010","111111111111011100","111111111111111100","111111111111111100","000000000000011101","111111111110110100","000000000000001000","000000000000011000","000000000000001100","000000000000001001","111111111111101000","000000000000101010","000000000000000000","000000000000001000","000000000000010111","111111111111111100","000000000000010101","111111111111100111","111111111111110010","000000000000100010","000000000000001001","111111111111111111","111111111111100101","111111111111110110","000000000000000001","000000000000000100","111111111111111000","000000000000000100","000000000000000010","111111111111101100","000000000000000000","111111111111011110","000000000000000001","000000000000010111","111111111111101111","000000000000001110","111111111111110110","000000000000010000","111111111111101110","000000000000011010","000000000000100011","000000000000000111","000000000000101111","111111111111010100","111111111111111001","111111111111101101","111111111111100001","111111111111111111","000000000000010000","000000000000011110","111111111111110100","111111111111100111","000000000000010110","000000000000000110","000000000000000000","000000000000000111","111111111111111011","000000000000001011","111111111111111101","111111111111011001","111111111111000010","111111111111011111","111111111111100101","000000000000000101","111111111111111000"),
("111111111111111000","000000000000011011","111111111110101111","000000000000010001","000000000000000001","000000000000010101","000000000000010011","111111111111100001","000000000000000000","111111111111110010","000000000000101101","111111111111101111","000000000000101101","111111111111010100","111111111111101100","000000000000001000","000000000000000101","000000000000100110","000000000000000101","000000000000011000","000000000000000100","000000000000011011","000000000000011110","111111111111111100","000000000000000111","000000000000011001","000000000000000110","000000000000000000","111111111111110011","000000000000011101","000000000000011011","000000000000000000","000000000000001001","111111111111110010","000000000000000000","111111111111111011","000000000000010110","111111111111111000","111111111111010111","000000000000010100","000000000000010100","111111111111111011","111111111110111000","111111111111011000","111111111111110111","111111111111110011","111111111111110000","111111111111101000","111111111111111001","111111111111101001","000000000000010011","000000000000011110","000000000000100000","111111111111111110","000000000000001111","111111111111100010","000000000000000011","000000000000001000","111111111111111001","111111111111111011","000000000000000111","111111111111111110","000000000000001001","111111111111111101","111111111111000101","111111111111110001","000000000000100100","111111111111111111","111111111110101101","000000000000000011","000000000000000101","000000000000010001","000000000000010100","000000000000000000","000000000000010100","111111111111111000","000000000000000011","111111111111111110","000000000000000011","000000000000001101","111111111111101010","000000000000000100","000000000000001010","111111111111111010","000000000000001001","111111111111010110","111111111111110111","000000000000010110","111111111111110001","000000000000001011","000000000000000001","111111111111111101","000000000000000011","000000000000000100","111111111111100101","111111111111011011","000000000000010000","000000000000000100","000000000000010000","000000000000001100","000000000000011010","111111111111111001","000000000000000001","000000000000011010","000000000000000111","000000000000011001","111111111111110000","111111111111101111","111111111111110001","111111111111110010","111111111111111111","000000000000001011","000000000000010100","000000000000000010","000000000000001000","000000000000000110","111111111111111010","000000000000011100","111111111111110111","000000000000001111","111111111111111110","000000000000001011","111111111111010100","111111111110111011","111111111111110101","111111111111110100","000000000000010111","000000000000000010"),
("111111111111101010","000000000000010100","111111111110101111","000000000000000110","111111111111100111","000000000000010101","000000000000100011","111111111111100000","000000000000000100","111111111111111011","000000000000011100","111111111111110000","000000000000101101","111111111111100001","111111111111000000","000000000000000100","111111111111111010","000000000000010000","000000000000000101","000000000000010001","111111111111101010","000000000000000101","000000000000000111","111111111111110010","111111111111111110","111111111111111101","000000000000100101","000000000000000010","111111111111110101","000000000000000000","111111111111110110","000000000000010001","000000000000000010","000000000000010011","000000000000011100","111111111111100011","111111111111111000","000000000000010100","111111111111101101","000000000000010101","000000000000010101","000000000000000101","111111111111001110","000000000000001011","000000000000000010","111111111111100001","111111111111101110","111111111111100110","000000000000000011","000000000000000011","000000000000000001","000000000000010001","000000000000010011","111111111111101010","000000000000001111","111111111111101010","000000000000000110","111111111111111100","111111111111111000","000000000000001111","000000000000001101","000000000000100111","000000000000001101","111111111111111101","111111111111010111","111111111111111110","000000000000011001","000000000000100000","111111111110111010","111111111111111010","111111111111111111","000000000000010100","000000000000010010","111111111111101010","000000000000100000","000000000000010010","000000000000000001","000000000000000111","111111111111111101","000000000000010001","000000000000001110","111111111111110010","111111111111111111","111111111111101101","111111111111111011","111111111111111001","111111111111011100","000000000000000001","111111111111101010","000000000000000110","111111111111110000","000000000000000100","111111111111101011","000000000000010011","111111111111110110","111111111111101000","000000000000010100","000000000000000001","000000000000100100","111111111111101100","000000000000010111","000000000000000100","000000000000000110","000000000000010001","000000000000010010","000000000000010001","111111111111001110","111111111111101101","111111111111011110","111111111111100000","111111111111111000","000000000000000100","000000000000000001","000000000000000000","111111111111100100","000000000000010110","000000000000011100","111111111111111100","111111111111011110","000000000000000001","000000000000001100","000000000000011001","111111111111101011","111111111111000000","111111111111110000","111111111111110110","000000000000001011","111111111111101111"),
("111111111111111011","000000000000001100","111111111110101010","111111111111110001","111111111111101110","000000000000010000","000000000000010101","000000000000001010","000000000000000011","000000000000001111","000000000000011011","000000000000001110","000000000000101001","111111111111111000","111111111110101111","111111111111111100","000000000000000101","000000000000010001","000000000000011111","111111111111111011","111111111111100111","000000000000010011","000000000000101011","000000000000000011","111111111111110011","000000000000010101","000000000000101000","111111111111111111","111111111111110010","111111111111101111","111111111111111010","111111111111101000","111111111111111011","000000000000011100","000000000000100110","111111111111110101","000000000000010111","000000000000001111","111111111111011000","111111111111100111","000000000000001001","000000000000100101","111111111111110011","000000000000101001","000000000000010010","111111111111010101","000000000000100101","000000000000000111","111111111111101110","000000000000000101","111111111111111010","000000000000000010","000000000000000011","111111111111100101","000000000000001100","111111111111010101","111111111111110000","000000000000001011","000000000000010110","000000000000000111","000000000000001100","000000000000100110","000000000000010101","111111111111101100","111111111111010101","000000000000010100","000000000000100000","000000000000011111","111111111110101001","000000000000000001","000000000000001101","111111111111101110","000000000000011001","111111111111110100","000000000000010100","000000000000001001","000000000000000011","000000000000000101","111111111111011101","000000000000000010","111111111111111010","000000000000000101","111111111111101111","111111111111111001","000000000000000110","111111111111011000","111111111111100011","000000000000100011","111111111111110000","111111111111111111","111111111111011000","111111111111101111","111111111111110110","000000000000011011","000000000000001101","111111111111110110","111111111111111111","111111111111111100","000000000000000010","000000000000000000","000000000000010010","000000000000100001","000000000000011101","111111111111101110","000000000000000110","000000000000100001","111111111111101110","000000000000001000","111111111111101010","111111111111101010","111111111111111000","000000000000010101","000000000000100010","111111111111111111","111111111111110111","000000000000010110","000000000000010100","000000000000000000","111111111111011010","000000000000001000","111111111111111001","000000000000101010","111111111111111011","111111111111101011","000000000000000111","000000000000010001","111111111111111101","111111111111101011"),
("000000000000000000","000000000000001011","111111111111010110","000000000000001001","111111111111111101","000000000000001110","111111111111101010","000000000000011111","111111111111100011","000000000000011001","000000000000100100","111111111111111100","000000000000000011","000000000000011010","111111111111100011","000000000000011110","000000000000000000","000000000000001001","000000000000010100","000000000000011001","111111111111110101","111111111111110000","000000000000111001","000000000000010000","111111111111110001","111111111111111101","000000000000011011","111111111111101011","111111111111010101","000000000000001111","000000000000001101","111111111111101111","000000000000010010","000000000000010001","000000000000010111","111111111111110011","000000000000011011","000000000000010111","111111111111011011","111111111111110011","000000000000001100","111111111111111100","000000000000011000","000000000000010110","111111111111110111","111111111111101110","000000000000011111","111111111111111000","111111111111110110","111111111111101111","111111111111101100","000000000000001000","000000000000001010","111111111111001101","000000000000101101","111111111111010101","111111111111101010","111111111111110010","111111111111111000","111111111111111101","111111111111110110","000000000000101001","000000000000001011","111111111111110110","111111111111100010","111111111111111111","000000000000001111","000000000000100001","111111111110100011","000000000000001101","111111111111111011","000000000000000101","000000000000100110","111111111111101001","000000000000000010","000000000000000111","000000000000001110","111111111111110100","111111111111101111","000000000000010101","111111111111111110","000000000000000001","111111111111100011","111111111111101100","000000000000010000","111111111111110010","111111111111101000","000000000000001010","000000000000000111","111111111111111111","111111111111111001","111111111111111101","000000000000001001","000000000000011100","000000000000001110","111111111111100101","000000000000001100","111111111111100110","000000000000001011","000000000000010000","000000000000010011","000000000000010111","111111111111101101","000000000000001010","000000000000000111","000000000000010110","111111111111010100","000000000000000001","111111111111101001","000000000000010001","111111111111100101","000000000000100011","000000000000100000","000000000000000110","111111111111001101","000000000000011011","000000000000000011","000000000000101000","111111111111100001","000000000000010011","000000000000000000","000000000000010110","000000000000010111","000000000000100110","000000000000000000","000000000000000100","000000000000011010","111111111111110101"),
("111111111111111100","000000000000000011","111111111111011100","000000000000000000","000000000000000000","000000000000011001","000000000000000010","000000000000100000","111111111111101011","000000000000101001","000000000000011100","111111111111111011","000000000000000100","000000000000011011","000000000000001100","000000000000010011","111111111111110110","000000000000001100","000000000000001001","000000000000000101","111111111111101100","111111111110110110","000000000000011111","000000000000001001","000000000000010010","000000000000000001","111111111111110101","111111111111111001","111111111111110010","000000000000010010","111111111111100110","111111111111110011","111111111111111011","000000000000010011","000000000000100011","111111111111011100","000000000000000110","000000000000000111","111111111111010000","111111111111101110","000000000000010101","111111111111111101","000000000000100000","000000000000001010","000000000000000100","000000000000001011","000000000000011010","111111111111110010","000000000000000000","111111111111101100","000000000000001110","000000000000001101","000000000000010010","111111111111001010","000000000000001010","111111111111110010","111111111111100110","111111111111110100","000000000000001110","111111111111110100","111111111111111101","000000000000011010","000000000000001101","111111111111101101","111111111111101110","000000000000001010","000000000000010101","000000000000000010","111111111110110101","000000000000001111","111111111111101000","111111111111111101","000000000000010001","111111111111100110","111111111111101010","000000000000001110","000000000000001100","000000000000001010","000000000000001000","000000000000000000","000000000000010110","111111111111111100","111111111111011101","000000000000001100","000000000000010100","000000000000001001","111111111111011000","000000000000101000","111111111111110001","111111111111110100","111111111111111000","111111111111111001","000000000000100001","000000000000011010","111111111111101011","111111111111101001","111111111111110000","111111111111110110","000000000000001010","000000000000011101","111111111111110001","000000000000101000","111111111111111100","000000000000001010","000000000000000110","000000000000000110","111111111111110001","111111111111111101","111111111111100100","111111111111110011","111111111111110010","000000000000010111","000000000000010011","111111111111100010","111111111111101000","000000000000000110","000000000000000110","000000000000010010","111111111111101111","000000000000011001","000000000000010011","000000000000000011","000000000000111001","000000000000100101","111111111111110000","000000000000011001","000000000000100000","111111111111111110"),
("111111111111110101","111111111111110101","000000000000010011","111111111111101101","111111111111100110","111111111111110001","000000000000000000","000000000000011000","111111111111111011","000000000000100110","000000000000010110","111111111111111000","000000000000000000","111111111111111001","111111111111111111","000000000000000111","000000000000001010","000000000000010001","000000000000001111","000000000000011000","000000000000001010","111111111110111001","000000000000000110","111111111111101000","000000000000010011","111111111111101100","111111111111110101","000000000000001101","000000000000000111","000000000000001000","000000000000000110","000000000000011001","000000000000011011","111111111111110110","000000000000000100","111111111111111000","111111111111111001","000000000000001110","111111111111011000","000000000000001001","111111111111111001","111111111111110111","000000000000010000","111111111111111111","111111111111110000","000000000000011011","000000000000000000","000000000000010110","000000000000000110","000000000000000001","000000000000001111","000000000000000001","111111111111101101","111111111111101111","000000000000000101","111111111111110011","111111111111111001","111111111111111100","111111111111111001","000000000000000011","000000000000001001","000000000000011010","000000000000001000","111111111111101000","111111111111111011","000000000000001101","000000000000100110","000000000000010101","111111111111010110","111111111111110010","000000000000001110","000000000000001111","000000000000100011","111111111111110110","000000000000000001","000000000000001010","111111111111111011","111111111111110111","111111111111110100","000000000000001000","111111111111111110","111111111111110010","111111111111101010","000000000000000100","000000000000000110","000000000000000011","111111111111011100","000000000000011100","111111111111111100","000000000000001111","000000000000000111","111111111111111000","000000000000011100","000000000000001011","111111111111110010","000000000000001000","000000000000010000","111111111111111011","000000000000000110","000000000000011101","111111111111101011","000000000000100100","000000000000010100","000000000000010010","111111111111111011","111111111111110111","111111111111011101","111111111111110101","111111111111011010","000000000000000000","000000000000000101","000000000000000110","000000000000001000","111111111111111001","000000000000000101","000000000000010001","000000000000011000","000000000000010101","000000000000000010","000000000000000100","000000000000011101","111111111111011010","000000000000010111","000000000000011000","111111111111101110","000000000000010001","111111111111111101","000000000000000110"),
("111111111111100111","000000000000000101","000000000000000100","000000000000010001","000000000000000101","000000000000001011","000000000000000011","000000000000010000","111111111111011011","000000000000000101","000000000000011101","111111111111011000","111111111111110101","111111111111001010","000000000000010010","000000000000010110","000000000000001100","111111111111111000","000000000000000111","111111111111111101","111111111111110101","111111111110100001","111111111111110101","111111111111100011","111111111111100011","111111111111110111","111111111111101101","111111111111110110","000000000000100011","000000000000011101","111111111111101000","000000000000001110","000000000000001101","000000000000000100","111111111111110000","111111111111100001","000000000000000000","000000000000001010","000000000000000010","000000000000001100","000000000000110001","000000000000000100","000000000000101111","000000000000000001","111111111111110101","000000000000010011","111111111111111110","000000000000000000","111111111111110000","000000000000001001","000000000000001010","000000000000000000","111111111111011100","111111111111111000","000000000000000011","111111111111100011","111111111111111111","000000000000000010","111111111111111001","000000000000001111","111111111111110011","000000000000001100","111111111111110111","111111111111100100","000000000000000000","000000000000001000","000000000000100101","000000000000001111","111111111111001100","111111111111101101","000000000000001100","000000000000000100","000000000000001110","000000000000010111","000000000000001101","000000000000011110","111111111111110011","111111111111111101","111111111111110111","000000000000001010","000000000000010100","111111111111110010","111111111111100101","000000000000001000","000000000000001110","000000000000011100","111111111111110000","000000000000010101","000000000000000010","000000000000000110","000000000000100101","111111111111111111","111111111111110110","000000000000010000","111111111111101010","000000000000000010","111111111111110100","111111111111110000","000000000000010101","000000000000001011","000000000000000010","111111111111111111","111111111111110011","000000000000000111","111111111111101101","111111111111111001","000000000000000111","111111111111111110","111111111111011011","111111111111110101","000000000000000001","000000000000010100","000000000000001010","000000000000000000","111111111111111101","000000000000011011","000000000000010100","000000000000100000","111111111111111000","000000000000010111","000000000000000000","111111111111110000","111111111111111101","000000000000011111","000000000000000000","000000000000001001","000000000000011000","000000000000010001"),
("111111111111101100","000000000000000000","111111111111110011","111111111111111100","000000000000001101","000000000000000000","111111111111100010","111111111111110111","111111111111100100","111111111111110010","000000000000001010","111111111111101000","000000000000011001","111111111111000000","000000000000010001","000000000000000000","000000000000000001","000000000000000011","000000000000000100","000000000000000111","000000000000000010","111111111111000100","000000000000000010","111111111111111010","111111111111101001","000000000000011101","111111111111101010","000000000000001000","000000000000001001","000000000000011010","000000000000000110","000000000000011000","000000000000000000","000000000000010101","000000000000001011","000000000000000101","000000000000000001","000000000000000111","000000000000001100","000000000000000000","000000000000010101","000000000000001000","000000000000011000","111111111111111101","111111111111111000","000000000000010011","000000000000010101","000000000000001101","000000000000001100","111111111111111010","111111111111110110","000000000000000010","111111111111011010","111111111111110111","111111111111110011","111111111111110000","000000000000010001","000000000000000000","111111111111111101","000000000000000010","000000000000000010","000000000000000000","000000000000000110","000000000000001001","111111111111100000","111111111111110111","000000000000010001","000000000000100111","000000000000001110","000000000000010000","000000000000011110","000000000000010111","111111111111101111","111111111111101110","000000000000010110","111111111111111111","000000000000000011","000000000000001000","111111111111110100","111111111111111010","000000000000010011","000000000000001010","111111111111110100","111111111111110000","111111111111111101","111111111111110010","000000000000011111","000000000000010110","111111111111110010","000000000000000000","000000000000100011","000000000000000110","000000000000011001","111111111111111101","111111111111101001","000000000000011000","000000000000000000","111111111111101011","000000000000011101","111111111111111101","111111111111111001","000000000000001010","000000000000010100","000000000000100010","111111111111010110","000000000000010010","111111111111101010","000000000000010010","111111111111110111","000000000000001000","111111111111111100","000000000000100101","000000000000001000","000000000000000001","000000000000010101","111111111111110011","000000000000010001","000000000000011110","111111111111110111","000000000000000011","000000000000010101","111111111111110111","000000000000000001","000000000000100110","111111111111101000","111111111111111000","111111111111111111","111111111111111010"),
("111111111111111000","000000000000000101","000000000000000010","000000000000001001","000000000000010000","000000000000000010","111111111111100001","111111111111011101","111111111111101010","000000000000010001","000000000000010111","111111111111101000","000000000000010101","111111111111001110","000000000000100011","000000000000011000","000000000000001110","111111111111111110","111111111111110110","000000000000010000","111111111111101000","000000000000010010","000000000000000000","111111111111101010","111111111111101101","000000000000000010","111111111111110001","111111111111111100","000000000000001010","000000000000011101","000000000000010100","000000000000010001","000000000000001001","000000000000010101","000000000000001011","000000000000000001","000000000000000101","000000000000101011","000000000000000000","111111111111111001","000000000000010100","111111111111101011","000000000000010001","111111111111111110","000000000000000000","111111111111111001","000000000000001101","000000000000001101","000000000000000010","000000000000001001","111111111111100111","000000000000001000","111111111111011111","111111111111111001","111111111111111111","000000000000001001","000000000000000000","000000000000000110","111111111111100110","000000000000001110","111111111111110010","000000000000010101","111111111111101010","111111111111100110","111111111111011100","111111111111110111","111111111111111010","111111111111111101","000000000000000100","111111111111110111","111111111111111010","000000000000001100","111111111111110000","000000000000001101","000000000000000011","111111111111110111","111111111111111010","000000000000001110","111111111111111110","000000000000000010","000000000000010110","111111111111111011","000000000000000100","111111111111101010","000000000000011111","000000000000000111","000000000000010001","000000000000001000","111111111111111010","111111111111111111","000000000000100001","000000000000000011","000000000000000010","111111111111111011","000000000000001000","111111111111111100","000000000000010010","111111111111101011","000000000000001101","111111111111110101","000000000000010011","111111111111111010","000000000000011011","000000000000011010","111111111111111001","111111111111100111","000000000000010011","000000000000001000","000000000000010011","111111111111100111","000000000000001000","000000000000101011","111111111111110001","000000000000001110","000000000000000011","111111111111110001","000000000000000010","000000000000001111","000000000000011011","000000000000010100","111111111111101111","000000000000000111","111111111111111101","000000000000011010","000000000000000100","000000000000000110","000000000000000110","000000000000000100"),
("000000000000011101","000000000000101100","000000000000100010","111111111111111111","111111111111111000","000000000000000000","111111111111110000","111111111111000010","111111111111111100","000000000000000000","000000000000100010","000000000000010001","000000000000010011","111111111111001101","000000000000001000","111111111111111101","000000000000000010","000000000000010001","000000000000000101","000000000000001001","111111111111110111","000000000000101110","000000000000100111","111111111111100011","000000000000000011","000000000000001010","111111111111110001","111111111111111010","111111111111111010","000000000000010011","000000000000100011","000000000000010101","111111111111110001","000000000000010011","000000000000000111","000000000000011110","111111111111101101","000000000000100000","000000000000000100","000000000000010011","000000000000010001","111111111111011011","000000000000010011","111111111111101110","000000000000000111","000000000000000001","111111111111111101","000000000000100000","111111111111110001","111111111111101000","111111111111100110","000000000000000110","111111111111101110","000000000000000010","000000000000001011","000000000000000010","000000000000010001","000000000000001010","111111111111101101","000000000000000110","000000000000011101","000000000000001101","000000000000000001","111111111111111101","111111111111011001","111111111111111010","111111111111111111","000000000000001010","111111111111101010","000000000000000011","000000000000011001","000000000000010001","111111111111100100","111111111111110001","000000000000010011","000000000000000110","000000000000000110","111111111111110100","111111111111101011","111111111111101011","000000000000011101","000000000000000001","111111111111111101","111111111111111001","000000000000101111","111111111111110000","111111111111111010","000000000000001001","111111111111111110","111111111111101001","000000000000011110","000000000000010010","000000000000010000","111111111111110010","111111111111110010","111111111111111000","111111111111110001","111111111111100010","111111111111111111","111111111111111110","111111111111110111","111111111111111100","000000000000100111","000000000000101101","111111111111100100","000000000000000010","000000000000000000","000000000000000100","000000000000000101","111111111111100001","000000000000001010","000000000000101001","000000000000001011","111111111111111100","000000000000100001","000000000000000011","111111111111111110","111111111111111011","000000000000000110","111111111111111110","000000000000001100","000000000000000011","111111111111101010","000000000000101010","000000000000000001","111111111111110000","111111111111111000","000000000000000111"),
("000000000000010111","000000000000101101","111111111111101000","000000000000001100","000000000000011100","000000000000011001","111111111111100000","111111111111101111","111111111111100001","111111111111111101","000000000000101000","000000000000000010","000000000000000011","111111111111011000","111111111111011011","111111111111111111","000000000000011110","000000000000100000","111111111111110110","000000000000001011","111111111111110101","000000000000001101","000000000000011010","111111111111110101","111111111111111111","000000000000000100","000000000000010001","111111111111111100","000000000000000101","000000000000011000","000000000000000010","000000000000000000","111111111111101100","000000000000101000","000000000000011000","000000000000011101","111111111111101101","000000000000001100","111111111111111111","000000000000010101","000000000000010101","111111111111101001","111111111111111010","000000000000010010","000000000000011010","000000000000001110","000000000000001001","000000000000001111","111111111111111100","000000000000000010","111111111111011010","000000000000000000","111111111111110010","000000000000100001","111111111111110111","111111111111110100","000000000000001101","111111111111100000","111111111111100010","000000000000010001","000000000000001111","111111111111110111","111111111111111011","000000000000000000","111111111111001011","111111111111110110","111111111111001101","000000000000011011","000000000000001111","000000000000000000","000000000000011000","000000000000000000","111111111111101110","000000000000001001","000000000000100000","000000000000000101","111111111111110011","111111111111110111","111111111111101001","111111111111011001","000000000000000000","000000000000010110","000000000000011000","111111111111011100","000000000000100110","111111111111110011","000000000000000001","000000000000000000","000000000000010001","000000000000011010","111111111111111111","111111111111111010","000000000000000000","111111111111111001","111111111111101100","111111111111100100","000000000000010010","111111111111110110","000000000000010110","111111111111110101","000000000000000011","000000000000000000","000000000000011011","000000000000011111","111111111111101110","111111111111111111","111111111111111101","111111111111111100","111111111111111001","111111111111101011","111111111111110100","000000000000100001","000000000000000011","111111111111111000","111111111111111000","111111111111110011","000000000000010110","000000000000000100","111111111111111100","000000000000000010","111111111111111010","000000000000000100","111111111111110010","000000000000010111","000000000000000010","111111111111111100","111111111111101000","000000000000010011"),
("000000000000101101","000000000000110100","000000000000000110","000000000000001100","111111111111100011","000000000000000101","111111111111110101","000000000000000111","000000000000001111","111111111111111100","000000000000001010","000000000000011000","000000000000000110","111111111111010111","111111111111110111","111111111111111011","000000000000000000","000000000000010000","000000000000010011","111111111111110100","000000000000000011","111111111111111001","000000000000011100","111111111111101110","000000000000000011","000000000000001110","111111111111110010","111111111111111011","111111111111110100","000000000000010001","000000000000011000","111111111111101110","111111111111101000","000000000000100100","000000000000010010","000000000000010110","111111111111101011","111111111111101010","000000000000001010","000000000000010110","000000000000000011","000000000000000100","000000000000010001","000000000000010001","111111111111111010","111111111111111001","111111111111111010","000000000000001101","111111111111111000","111111111111110100","111111111111101101","111111111111101110","111111111111110001","000000000000100101","000000000000000011","111111111111111111","000000000000000011","111111111111110010","111111111111110000","111111111111101110","000000000000000010","000000000000011100","000000000000001100","000000000000000101","111111111111011100","000000000000000000","111111111110001011","111111111111111011","000000000000010100","000000000000001110","000000000000100100","000000000000100001","111111111111011110","000000000000000011","000000000000100100","111111111111111010","000000000000000101","111111111111111010","111111111111101110","111111111111100011","111111111111110001","111111111111101110","000000000000001011","111111111111010101","000000000000100010","111111111111101001","000000000000000110","000000000000001010","111111111111111001","111111111111111101","000000000000001111","000000000000011000","111111111111100001","000000000000000101","111111111111110001","111111111111010101","000000000000000101","111111111111111000","111111111111101010","111111111111111101","000000000000010011","000000000000000110","111111111111110001","000000000000010011","111111111111110101","111111111111111111","000000000000000001","111111111111011010","111111111111111010","111111111111111100","111111111111110000","000000000000011011","000000000000010110","111111111111111000","111111111111110111","000000000000000100","111111111111101100","111111111111111010","111111111111110100","000000000000001111","000000000000010101","111111111111111101","111111111111101011","000000000000100001","111111111111011101","000000000000000000","111111111111101110","000000000000000111"),
("000000000000010110","000000000000010110","000000000000000010","111111111111111111","000000000000001010","000000000000010001","111111111111100110","000000000000001010","000000000000010000","111111111111111011","000000000000000001","000000000000101001","000000000000000011","111111111111110101","111111111111001010","111111111111110010","000000000000000110","000000000000001100","111111111111111110","000000000000011001","000000000000000111","111111111111100101","000000000000011000","111111111111110001","111111111111111000","000000000000000110","111111111111110001","000000000000000011","000000000000010110","111111111111111110","000000000000001111","000000000000000001","000000000000000000","111111111111110111","111111111111110000","000000000000011110","111111111111100110","000000000000010111","000000000000000100","000000000000000101","000000000000000011","111111111111101101","111111111111110101","000000000000010001","000000000000010101","111111111111100100","000000000000000100","000000000000101011","000000000000001010","111111111111111110","111111111111110000","000000000000001000","111111111111110101","000000000000011000","000000000000011001","111111111111101101","111111111111011001","111111111111100001","111111111111101110","111111111111110111","111111111111011000","000000000000001001","000000000000001010","111111111111110110","111111111111101000","111111111111101111","111111111110010110","111111111111110101","000000000000010011","111111111111110100","000000000000011100","000000000000001101","111111111111000100","000000000000000101","000000000000100111","000000000000000101","111111111111111101","111111111111110010","111111111111011011","000000000000000001","111111111111110110","111111111111111110","000000000000001000","111111111111000100","000000000000100100","111111111111010101","111111111111101100","111111111111110111","000000000000010000","000000000000000011","111111111111111000","000000000000001011","111111111111100100","000000000000011011","000000000000001101","111111111111011100","000000000000001100","111111111111101100","000000000000000000","111111111111111000","000000000000001001","111111111111111000","111111111111110101","000000000000011000","111111111111101101","111111111111111011","111111111111101000","111111111111001000","111111111111101100","111111111111100101","111111111111111100","000000000000000100","000000000000010010","000000000000000110","111111111111101001","111111111111110100","000000000000000001","111111111111101011","111111111111001000","000000000000000100","111111111111111101","000000000000000001","111111111111101010","000000000000001110","111111111111101011","111111111111111111","111111111111110110","111111111111111100"),
("000000000000011101","000000000000000110","111111111111111001","000000000000000110","000000000000010010","000000000000100111","111111111111110111","000000000000100010","000000000000010010","111111111111110000","000000000000000001","000000000000100110","000000000000000100","111111111111111011","111111111111010111","111111111111111100","000000000000001100","000000000000010100","111111111111110110","000000000000000100","111111111111100111","111111111111110101","000000000000011001","111111111111011100","111111111111101001","000000000000100010","111111111111111011","111111111111111110","000000000000001111","111111111111101100","000000000000000100","111111111111110010","000000000000000101","000000000000001111","000000000000000110","000000000000001010","111111111111111011","111111111111111011","111111111111111001","111111111111111111","111111111111110111","111111111111101010","000000000000000000","111111111111111001","000000000000001011","111111111111111001","111111111111001111","000000000000010110","000000000000000000","111111111111011101","000000000000000001","000000000000000111","000000000000000000","000000000000001111","111111111111111011","111111111111110011","111111111111011010","111111111111110001","000000000000000101","111111111111110111","111111111111000101","000000000000001001","111111111111110100","000000000000001101","000000000000010101","111111111111111000","111111111110111011","000000000000000000","000000000000010001","111111111111101101","000000000000010010","000000000000011010","111111111110111110","111111111111111101","000000000000100010","000000000000000101","111111111111111110","111111111111110001","111111111111011000","000000000000011000","111111111111100011","000000000000001010","111111111111111010","111111111111101111","000000000000011000","111111111111011010","111111111111101010","000000000000001100","000000000000010100","000000000000010001","000000000000001100","111111111111111001","000000000000001000","000000000000001110","111111111111111101","111111111111000010","111111111111011010","111111111111110000","111111111111001010","000000000000000101","000000000000011000","000000000000000000","111111111111011110","000000000000001001","111111111111110110","000000000000010001","111111111111111001","111111111111010100","111111111111101100","111111111111011011","111111111111110011","000000000000001110","000000000000000111","000000000000001000","000000000000011000","111111111111110011","111111111111100100","000000000000001000","111111111111000010","000000000000011001","000000000000010111","111111111111111100","111111111111111000","000000000000010110","111111111111101000","000000000000001100","111111111111111000","000000000000000111"),
("000000000000101001","000000000000100001","111111111111100100","000000000000010111","111111111111111000","000000000000011011","111111111111111110","000000000000011100","111111111111111101","000000000000001001","111111111111110011","000000000000001100","000000000000100100","000000000000000111","111111111110111001","000000000000001011","111111111111111100","000000000000011110","111111111111011001","000000000000010011","000000000000001011","000000000000000010","000000000000000100","111111111111011110","000000000000000000","000000000000011101","000000000000011011","000000000000001100","111111111111101110","111111111111100110","111111111111111100","111111111111011000","111111111111100100","000000000000010110","111111111111111110","111111111111110001","111111111111110100","000000000000001101","000000000000000011","111111111111101010","000000000000100100","000000000000000000","111111111111110000","000000000000001011","000000000000000100","111111111111100000","111111111111100101","000000000000100000","000000000000000000","111111111111110110","000000000000010101","000000000000001111","111111111111100011","000000000000011001","000000000000010011","000000000000000000","111111111111011101","111111111111010011","111111111111110101","111111111111110111","111111111110111010","111111111111101111","000000000000010010","000000000000000111","000000000000001001","111111111111110010","111111111111011110","111111111111110101","111111111111110010","111111111111101000","000000000000100100","111111111111110110","111111111111001001","000000000000001011","000000000000011100","111111111111111100","000000000000010001","111111111111101001","111111111111001010","111111111111100111","111111111111111010","000000000000001010","111111111111111010","111111111111101111","000000000000011101","111111111111010010","000000000000000110","000000000000010001","000000000000010111","111111111111100110","111111111111100101","111111111111110110","111111111111101100","000000000000001110","111111111111110000","111111111111110100","111111111111111101","000000000000001010","111111111111010010","111111111111110001","000000000000100000","000000000000000000","111111111111010010","000000000000011100","111111111111100110","000000000000000011","111111111111110111","111111111111100111","111111111111101111","111111111111010101","000000000000000010","000000000000001100","000000000000010000","111111111111111101","111111111111111111","000000000000000011","111111111111011010","111111111111111111","111111111111101100","000000000000001111","000000000000011010","000000000000001111","111111111111011101","111111111111101110","111111111111100100","000000000000010100","111111111111111000","111111111111101110"),
("000000000000100110","000000000000010010","000000000000010101","000000000000011111","111111111111101110","000000000000001110","000000000000000011","000000000000011011","000000000000100001","111111111111111101","000000000000010001","000000000000000101","000000000000011101","000000000000010001","111111111111100100","111111111111111111","111111111111011100","000000000000000110","111111111111111101","111111111111111101","000000000000000100","111111111111010001","111111111111111100","111111111111110011","000000000000000000","000000000000110011","000000000000100000","000000000000010000","000000000000000011","111111111111010011","000000000000011100","111111111111110010","000000000000000001","111111111111111011","000000000000001101","000000000000000111","111111111111111111","000000000000000110","111111111111101110","111111111111111011","000000000000001011","111111111111100111","111111111111111100","111111111111111000","000000000000000000","111111111111110011","111111111111100011","111111111111111101","111111111111011011","111111111111100101","111111111111110010","111111111111101101","111111111111100100","000000000000101010","000000000000001100","000000000000001111","111111111111011000","111111111111111110","111111111111010111","111111111111111111","111111111111011101","000000000000000011","000000000000010011","111111111111111111","000000000000011010","111111111111011011","111111111111011000","111111111111011111","111111111111110100","111111111111101101","000000000000010010","000000000000001100","111111111111011011","111111111111111000","000000000000001011","000000000000000010","000000000000000100","111111111111101101","111111111111011100","111111111111111110","111111111111100110","111111111111111101","111111111111111000","111111111111100110","000000000000100001","111111111111110100","000000000000000010","000000000000100100","000000000000011000","111111111111110010","000000000000001010","111111111111101101","111111111111101110","111111111111101111","111111111111111001","111111111111101001","000000000000010110","000000000000001000","111111111111010100","111111111111110100","000000000000010110","111111111111111111","111111111111000111","000000000000000101","111111111111100011","000000000000001110","111111111111111011","111111111111110100","111111111111100110","111111111111010111","111111111111111110","111111111111110010","000000000000000011","111111111111101000","000000000000011011","111111111111111110","111111111111011010","111111111111111000","111111111111101101","111111111111111010","000000000000000010","111111111111111110","111111111111101000","000000000000001100","111111111111110011","111111111111111000","111111111111101011","111111111111110000"),
("000000000001001101","000000000000010110","000000000000001110","111111111111111010","111111111111111000","111111111111111111","000000000000001011","111111111111011111","111111111111110111","111111111111110000","111111111111111010","111111111111101100","000000000000100011","000000000000100111","000000000000001001","111111111111110100","111111111111111100","000000000000001001","111111111111100101","111111111111101100","000000000000111000","111111111111001100","111111111111101101","000000000000001111","000000000000000011","000000000000000100","111111111111101100","000000000000000000","000000000000000111","111111111111011111","000000000000001101","111111111111110011","111111111111111001","000000000000010011","111111111111111010","000000000000000000","000000000000001101","111111111111111101","111111111111010111","111111111111101011","000000000000011111","111111111111011110","111111111111111110","000000000000010011","111111111111110001","000000000000000100","111111111111010011","000000000000010111","111111111111010001","111111111111110101","111111111111111110","111111111111111110","111111111111111111","000000000001000100","000000000000001101","000000000000010011","111111111111100010","111111111111111110","111111111111100110","111111111111111001","111111111111100010","000000000000000011","000000000000010001","111111111111111110","000000000000101001","111111111111100100","000000000000000000","111111111111100110","111111111111110100","111111111111010111","000000000000010100","000000000000000111","000000000000001111","000000000000001001","111111111111111001","000000000000000010","111111111111111110","111111111111111000","111111111111110110","111111111111111000","111111111111101111","000000000000000000","000000000000010100","111111111111001010","000000000000011100","111111111111100111","111111111111111101","000000000000011001","111111111111101111","111111111111101000","000000000000010110","111111111111110000","111111111111100010","000000000000000100","000000000000100100","000000000000010000","000000000000100011","000000000000001100","000000000000000111","111111111111111000","111111111111110100","111111111111101000","111111111111101000","111111111111111111","000000000000000000","111111111111111110","000000000000000011","000000000000000001","111111111111001101","111111111111110000","000000000000000101","000000000000001000","111111111111011110","111111111111101101","111111111111100111","111111111111111011","111111111111101010","111111111111100111","111111111111010010","111111111111011110","111111111111111110","000000000000000000","000000000000011111","000000000000101011","000000000000010100","000000000000100101","111111111111100101","111111111111100011"),
("000000000000100101","000000000000100010","000000000000100010","111111111111110111","000000000000000010","111111111111111011","111111111111111110","111111111111110001","111111111111110111","111111111111100001","000000000000011010","000000000000000011","000000000000011010","000000000000111000","111111111111100010","000000000000000001","000000000000000010","000000000000101000","000000000000000100","111111111111111000","000000000000110110","111111111111010010","111111111111101100","000000000000000000","000000000000001010","000000000000100000","111111111111100100","111111111111110001","000000000000001010","111111111111101100","000000000000111101","000000000000001011","111111111111100001","111111111111110100","000000000000010001","111111111111111011","000000000000010010","000000000000011101","111111111111100011","111111111111100100","111111111111011110","111111111111110001","111111111111111010","000000000000001011","111111111111010111","000000000000010101","111111111111011010","000000000000001001","111111111111001101","111111111111011100","111111111111001110","111111111111011101","111111111111110110","000000000000101100","111111111111111100","111111111111100110","000000000000000000","111111111111110100","111111111111000000","000000000000001010","111111111111111100","000000000000001000","000000000000000010","000000000000000000","000000000000001111","111111111111111000","000000000000001011","111111111111111111","000000000000000001","111111111111100100","000000000000001010","000000000000000110","000000000000001011","111111111111111101","000000000000010011","111111111111100001","111111111111111100","111111111111110001","111111111111010111","111111111111100001","000000000000011101","111111111111111111","000000000000000111","111111111111001000","000000000000011001","111111111111100011","000000000000001011","000000000000010011","000000000000000000","111111111111110101","111111111111101001","111111111111100010","000000000000011101","000000000000001010","111111111111011010","000000000000010010","111111111111110001","000000000000100000","000000000000000011","111111111111101001","000000000000001010","000000000000001101","111111111111111101","000000000000000101","000000000000000011","111111111111110011","000000000000000111","111111111111111011","111111111111110101","111111111111010110","000000000000000011","000000000000110001","111111111111111010","111111111111100101","111111111111011001","111111111111111110","111111111111110010","000000000000001100","000000000000000000","111111111111100100","000000000000001101","000000000000011001","000000000000000110","000000000000000100","111111111111111111","000000000000101110","000000000000001000","111111111111111110"),
("111111111111110001","111111111111010010","111111111111101000","000000000000001001","000000000000010000","000000000000101110","111111111111111101","000000000000011111","000000000000010010","000000000000000000","000000000000011010","111111111111100011","000000000000011001","111111111111111111","111111111111101001","111111111111110111","000000000000100011","000000000000001010","111111111111011001","000000000000000000","111111111111111011","111111111111101100","000000000000010110","000000000000000000","111111111111110010","000000000000001100","000000000000000100","000000000000000000","000000000000010100","000000000000010010","000000000000000111","000000000000001000","111111111111101101","111111111111110010","000000000000000110","000000000000011001","000000000000000010","000000000000010101","111111111111100011","111111111111110111","111111111111101000","000000000000000101","000000000000001111","000000000000100011","111111111111111110","000000000000011110","111111111111100100","000000000000010111","111111111111101110","111111111111100100","111111111111110110","000000000000000000","111111111111110001","000000000000000000","000000000000011100","000000000000000001","000000000000001001","111111111111110001","111111111111110100","000000000000000000","111111111111110101","000000000000000111","000000000000011011","000000000000010010","000000000000100010","111111111111011101","000000000000100101","111111111111110101","000000000000001100","111111111111101010","000000000000100010","000000000000100000","000000000000000101","000000000000001001","111111111111111100","000000000000001101","111111111111111101","111111111111111110","000000000000000011","111111111111110001","000000000000000000","111111111111101010","000000000000001111","000000000000000000","000000000000011100","111111111111110110","111111111111111011","000000000000001101","111111111111011110","000000000000000100","000000000000000000","111111111111100010","111111111111101100","000000000000011101","111111111111010101","111111111111101010","111111111111100101","111111111111101111","000000000000011111","000000000000000111","111111111111110001","000000000000000000","111111111111100001","111111111111101100","111111111111111000","000000000000000000","000000000000001000","000000000000000101","000000000000000000","111111111111111101","111111111111101001","000000000000010110","111111111111111111","111111111111110100","000000000000001000","111111111111110010","111111111111111110","000000000000000101","000000000000001011","111111111111110111","111111111111110110","000000000000010000","111111111111110111","000000000000100010","000000000000010011","111111111111111000","000000000000000011","000000000000011000"),
("000000000000000010","000000000000010010","000000000000001000","000000000000010001","000000000000001111","111111111111111011","111111111111110001","000000000000010000","111111111111110110","111111111111111110","000000000000000110","000000000000000111","000000000000000100","111111111111111100","000000000000001001","111111111111110101","111111111111111101","000000000000001010","111111111111110001","111111111111110011","000000000000000000","000000000000001011","000000000000000000","111111111111110000","111111111111110011","000000000000000000","000000000000000101","000000000000000111","111111111111111000","000000000000000011","111111111111111010","111111111111111010","111111111111111101","000000000000000111","000000000000000011","000000000000010101","000000000000001100","000000000000001110","000000000000010000","000000000000010010","000000000000001111","000000000000001111","000000000000010001","000000000000011000","111111111111101111","111111111111110100","000000000000010000","000000000000001011","000000000000000111","111111111111110100","000000000000001011","111111111111100111","111111111111101011","111111111111110101","000000000000000111","111111111111110101","000000000000010100","111111111111111000","000000000000001010","111111111111110111","000000000000001011","000000000000001110","111111111111101011","111111111111101111","000000000000011000","000000000000000011","000000000000001001","000000000000000000","000000000000010000","000000000000001011","111111111111111000","000000000000010010","111111111111111010","111111111111101111","000000000000000101","111111111111101111","111111111111101110","111111111111111110","111111111111111010","111111111111101001","111111111111111010","111111111111101010","000000000000010000","111111111111111111","000000000000010010","000000000000010100","000000000000001100","111111111111110100","000000000000000001","000000000000001100","000000000000010000","111111111111101110","111111111111101011","111111111111111110","111111111111111110","000000000000000111","000000000000000101","000000000000001101","000000000000000001","000000000000000100","000000000000000011","111111111111111100","000000000000000100","111111111111110101","000000000000000000","111111111111101101","000000000000000010","111111111111111010","111111111111110100","000000000000000111","111111111111110100","111111111111111110","111111111111111001","111111111111101011","000000000000000110","111111111111101011","000000000000000110","000000000000001101","000000000000000110","111111111111111100","111111111111110001","000000000000010110","000000000000001001","111111111111111011","111111111111110011","111111111111111000","000000000000000011","000000000000000010"),
("111111111111111011","000000000000001110","000000000000001101","111111111111110100","111111111111110110","111111111111111110","111111111111111101","000000000000001111","000000000000010000","000000000000000010","000000000000000001","111111111111101101","111111111111110100","000000000000000111","111111111111101011","111111111111111001","111111111111110101","000000000000010101","111111111111101011","111111111111111100","111111111111111110","000000000000001011","000000000000010011","111111111111110110","000000000000000001","000000000000001101","111111111111110011","111111111111110100","000000000000010001","000000000000010111","000000000000001100","000000000000010100","111111111111101100","000000000000001101","000000000000010100","111111111111110100","111111111111111001","000000000000001011","111111111111110110","000000000000000010","111111111111110111","111111111111111001","000000000000010011","000000000000001001","111111111111101000","111111111111111011","000000000000010100","111111111111110010","111111111111100111","000000000000001100","000000000000001101","000000000000000000","111111111111110110","000000000000000000","111111111111110110","000000000000001001","111111111111110111","111111111111100110","000000000000001011","000000000000001111","000000000000001011","000000000000010011","000000000000010001","000000000000010011","111111111111111001","000000000000000101","111111111111110000","111111111111110000","111111111111111011","111111111111110110","000000000000000000","000000000000010010","000000000000000000","111111111111110001","000000000000010111","000000000000001011","000000000000001011","000000000000000001","000000000000001000","111111111111110011","000000000000000101","000000000000000110","111111111111110000","000000000000001111","111111111111110101","111111111111110011","111111111111111101","000000000000001110","111111111111111010","000000000000011000","000000000000000000","000000000000001001","111111111111101101","000000000000011010","111111111111100110","111111111111110011","000000000000010010","000000000000000001","111111111111110100","000000000000001100","111111111111101011","111111111111111101","000000000000001011","111111111111110101","000000000000010101","000000000000000100","000000000000010001","111111111111111110","000000000000010111","000000000000000000","000000000000000100","111111111111110110","111111111111101010","111111111111110010","000000000000000100","000000000000000100","111111111111111100","111111111111111100","000000000000000000","111111111111111001","111111111111101011","000000000000010101","111111111111110110","111111111111110001","111111111111110101","111111111111110101","111111111111111001","111111111111110011"),
("000000000000001111","111111111111101110","000000000000001101","000000000000010000","111111111111111100","111111111111110111","111111111111110111","000000000000010011","000000000000011100","000000000000010100","000000000000001001","111111111111110110","000000000000000000","000000000000010001","000000000000001011","000000000000001010","111111111111111010","111111111111111000","000000000000000010","111111111111111110","111111111111111100","000000000000000000","000000000000011101","111111111111011111","111111111111111010","000000000000011010","000000000000000011","000000000000001010","000000000000010101","111111111111101011","000000000000001010","000000000000010101","111111111111110001","111111111111011011","000000000000001101","111111111111111001","000000000000001100","111111111111110001","000000000000000110","000000000000001010","111111111111111111","000000000000001100","111111111111110110","111111111111111000","000000000000000011","000000000000001110","000000000000001101","111111111111101011","111111111111101101","000000000000000101","000000000000000101","111111111111101111","111111111111111100","111111111111111010","000000000000000000","000000000000001000","111111111111011100","000000000000001000","000000000000001111","111111111111101111","000000000000010000","000000000000100000","000000000000010100","111111111111111100","111111111111110101","111111111111110001","111111111111110111","000000000000001100","000000000000010110","000000000000001010","000000000000010010","000000000000001111","111111111111011110","000000000000010011","111111111111101111","000000000000001100","111111111111111001","000000000000010100","111111111111110111","000000000000010111","111111111111100111","000000000000000001","000000000000010100","000000000000001010","000000000000000011","111111111111101010","111111111111100100","000000000000001111","111111111111111000","111111111111111010","000000000000001100","000000000000010001","000000000000000001","000000000000000101","111111111111101110","000000000000001001","000000000000011011","000000000000011110","111111111111110101","000000000000000110","111111111111110010","000000000000000110","000000000000001101","000000000000010000","111111111111101000","000000000000010100","000000000000001100","111111111111101111","000000000000000010","111111111111111111","000000000000000000","000000000000000000","111111111111110110","000000000000010011","000000000000000101","000000000000000100","000000000000010000","111111111111111110","000000000000001101","000000000000000101","111111111111100111","111111111111110111","111111111111110010","111111111111110110","000000000000011000","111111111111110001","000000000000000001","111111111111110010"),
("111111111111110111","111111111111110111","111111111111110001","000000000000100000","111111111111110001","000000000000001110","000000000000001101","000000000000010010","000000000000101000","111111111111011111","000000000000100111","111111111111111110","000000000000010000","111111111111011010","000000000000000000","000000000000010001","000000000000110100","000000000000000000","000000000000011110","000000000000110101","111111111111101101","111111111111111011","000000000000001110","111111111111111011","111111111111011000","000000000000010000","111111111111110111","000000000000110101","000000000000001011","111111111111100111","000000000000001001","111111111111101011","000000000000001001","111111111111101011","000000000000001001","111111111111111111","111111111111110011","000000000000010101","000000000000001111","111111111111100000","111111111111101001","111111111111010010","111111111111111111","111111111111111010","000000000000001000","000000000000000001","000000000000010010","111111111111101101","111111111111101101","111111111111101000","000000000000000110","000000000000100000","111111111111100100","000000000000000010","000000000000010011","000000000000000111","111111111111110000","000000000000000110","111111111111011111","000000000000001010","111111111111011101","000000000000011110","000000000000010101","000000000000000000","000000000000001000","111111111111110011","111111111111110001","000000000000000001","000000000000000100","111111111111111100","000000000000001100","000000000000000010","111111111111110111","000000000000000000","111111111111101000","000000000000001001","111111111111111100","000000000000100010","000000000000001110","000000000000101111","000000000000000110","000000000000001111","000000000000100100","111111111111101111","000000000000010100","111111111111011000","111111111111110110","111111111111111000","000000000000010101","111111111111110111","000000000000001110","111111111111110011","111111111111101001","000000000000001100","111111111111001011","000000000000001110","000000000000000110","000000000000000000","111111111111010100","111111111111011011","000000000000000010","000000000000001100","000000000000001010","000000000000000000","111111111111111100","000000000000001101","111111111111101110","111111111111010100","000000000000001110","000000000000001011","111111111111101000","000000000000011101","000000000000001100","111111111111111000","000000000000011111","000000000000100011","000000000000000010","000000000000000101","000000000000010010","111111111111110110","000000000000101010","000000000000001100","111111111111110010","111111111111110111","000000000000011001","111111111111111101","000000000000010111","111111111111011101"),
("111111111111100101","111111111111010110","111111111111011100","000000000000101011","000000000000010100","000000000000100101","111111111111111011","000000000000010000","000000000000100111","111111111111011010","000000000000100111","111111111111110001","000000000000010001","111111111111101001","111111111111101001","000000000000010111","000000000001000010","000000000000011011","000000000000011110","000000000000100010","111111111111011010","000000000000000000","000000000000010010","111111111111010001","111111111111101010","000000000000010111","111111111111011100","000000000000100000","000000000000010011","000000000000000001","000000000000000000","111111111111110110","000000000000001100","000000000000000011","111111111111101100","111111111111111100","111111111111011000","000000000000011111","000000000000000010","111111111111110001","000000000000000110","000000000000001000","111111111111101011","111111111111100100","000000000000010101","111111111111110100","000000000000110000","111111111111101110","111111111111110110","111111111111110001","000000000000010011","000000000000011100","111111111111100110","000000000000000011","000000000000011001","111111111111110001","111111111111110010","000000000000001011","111111111111100101","111111111111111101","111111111111111011","000000000000100101","000000000000111000","000000000000010001","111111111111111011","111111111111101110","111111111111011111","000000000000001001","000000000000000111","111111111111101011","000000000000100000","000000000000001110","111111111111011010","000000000000000011","000000000000001001","000000000000000001","000000000000000100","000000000000101101","111111111111011000","000000000000011011","000000000000001001","000000000000011000","000000000000110011","000000000000000010","000000000000110000","111111111111111110","111111111111110111","000000000000000000","111111111111100110","111111111111111001","111111111111100001","111111111111111001","111111111111101111","000000000000000010","111111111111101011","000000000000000110","000000000000001000","000000000000001100","111111111111110011","111111111111011011","000000000000001001","000000000000000101","000000000000010110","000000000000101111","111111111111010010","000000000000011000","111111111111011110","111111111111110100","000000000000101000","111111111111111100","111111111111011010","000000000000001011","111111111111110100","111111111111110000","111111111111111110","000000000000100111","000000000000000100","111111111111111011","111111111111111110","000000000000001010","000000000000010000","000000000000010011","000000000000000010","111111111111001001","000000000000001000","111111111111111101","000000000000001001","000000000000000000"),
("000000000000010000","111111111111100000","111111111111010110","000000000000001011","000000000000011111","000000000000000010","111111111111011101","000000000000000000","000000000000010001","111111111111110000","000000000000100000","000000000000001000","000000000000011100","111111111111101110","111111111111100001","000000000000000011","111111111111111011","000000000000001111","000000000000000000","000000000000000010","000000000000001010","111111111111110100","000000000000010001","111111111111001001","111111111111101111","111111111111111011","111111111111011000","111111111111111010","000000000000000000","000000000000010100","000000000000011110","111111111111111001","000000000000000110","000000000000011011","111111111111101011","000000000000000101","000000000000000101","000000000000001011","000000000000010010","000000000000000101","000000000000011101","000000000000010110","111111111111111011","111111111111100100","000000000000000111","111111111111100000","000000000000000001","111111111111111001","000000000000000011","111111111111111011","111111111111101111","000000000000011111","000000000000000000","000000000000000011","000000000000001000","111111111111111010","111111111111111111","000000000000001101","111111111111110110","111111111111111111","111111111111110000","111111111111111001","111111111111110110","111111111111100111","000000000000010000","111111111111110011","111111111111111010","000000000000010011","111111111111111001","111111111111111010","000000000000011010","111111111111111111","111111111111100101","111111111111110010","000000000000010011","111111111111111001","000000000000001010","000000000000010100","111111111111111011","111111111111110111","111111111111110100","000000000000000111","000000000000001000","000000000000010010","000000000000010011","111111111111110100","111111111111101011","000000000000000110","111111111111110011","111111111111101100","000000000000001111","111111111111111000","111111111111000000","000000000000010010","111111111111100111","000000000000011100","111111111111110100","000000000000010101","111111111111100101","111111111111100110","000000000000001110","111111111111101101","000000000000000000","000000000000000101","111111111111011101","111111111111111101","000000000000000000","111111111111110111","000000000000100001","000000000000001011","111111111111110011","000000000000010100","111111111111101100","000000000000000010","000000000000010100","000000000000000000","111111111111100111","000000000000000001","111111111111111001","000000000000011000","000000000000000001","000000000000011100","000000000000000000","111111111110110101","000000000000001001","111111111111111100","111111111111110000","000000000000010001"),
("000000000000001000","111111111111101011","111111111111000111","000000000000001101","000000000000010010","000000000000001000","000000000000000110","111111111111111101","000000000000010011","111111111111110011","000000000000011100","111111111111101011","000000000000011010","111111111111110100","111111111111111001","111111111111110011","111111111111110001","000000000000010000","111111111111101110","000000000000001001","000000000000001100","000000000000011110","000000000000001101","111111111111101010","000000000000001111","111111111111111001","111111111111110011","000000000000000011","111111111111110011","000000000000000111","000000000000101001","000000000000000000","000000000000000010","111111111111111011","000000000000000001","000000000000011101","000000000000000100","111111111111111001","000000000000011011","111111111111111010","000000000000011010","000000000000000111","111111111111011101","111111111110110101","000000000000000111","000000000000000101","111111111111011111","111111111111101101","111111111111100110","000000000000000100","000000000000001101","000000000000000110","111111111111111011","000000000000010010","111111111111110001","000000000000001101","000000000000010101","000000000000001001","111111111111111101","111111111111101110","111111111111101110","000000000000000011","000000000000000101","000000000000000010","111111111111010110","000000000000000101","000000000000001000","111111111111011010","000000000000001000","111111111111100111","111111111111110010","000000000000000000","111111111111100011","111111111111100000","000000000000011001","111111111111111010","111111111111111011","111111111111101110","111111111111111010","000000000000000100","000000000000000011","000000000000000010","111111111111111110","000000000000011001","000000000000001110","111111111111100001","111111111111111011","111111111111111011","111111111111111111","111111111111111100","111111111111110001","111111111111110000","111111111111110011","111111111111110110","111111111111101101","000000000000010111","111111111111111010","111111111111110000","111111111111111100","111111111111011011","111111111111101111","111111111111111010","111111111111100101","000000000000010010","111111111111100101","000000000000000111","000000000000010001","111111111111111011","000000000000101110","000000000000010101","000000000000000011","000000000000001100","111111111111011011","111111111111100001","111111111111111001","111111111111110010","111111111111011101","000000000000001110","000000000000001100","000000000000000001","111111111111110100","000000000000001010","111111111111010110","111111111110111010","111111111111101111","111111111111111011","000000000000010011","000000000000010101"),
("111111111111110100","111111111111111010","111111111111001111","000000000000000100","000000000000011100","111111111111101101","000000000000001111","000000000000000111","000000000000001010","111111111111111011","000000000000000110","111111111111110001","111111111111111010","111111111111001011","111111111111110111","111111111111110110","111111111111011010","000000000000001001","000000000000000011","000000000000000111","000000000000010001","000000000000110110","000000000000010001","111111111111110011","111111111111110110","000000000000010011","111111111111101110","000000000000001101","111111111111110010","111111111111110111","000000000000011010","000000000000011000","000000000000001001","000000000000000111","000000000000001101","000000000000000110","111111111111111100","000000000000010101","000000000000001001","000000000000001000","000000000000011110","111111111111110011","111111111111000010","111111111111010000","000000000000000110","111111111111101100","111111111111101000","111111111111110011","000000000000001001","000000000000000111","000000000000011011","000000000000010000","111111111111111111","000000000000010101","000000000000010011","111111111111101011","000000000000011100","111111111111101111","000000000000001001","111111111111110010","000000000000010111","111111111111110011","111111111111110101","000000000000010110","111111111110111110","111111111111101100","000000000000011001","111111111111101000","111111111111111111","111111111111111110","000000000000001101","000000000000001011","111111111111100111","111111111111010111","000000000000011001","000000000000000010","000000000000010001","111111111111110110","111111111111100010","111111111111110001","111111111111100101","000000000000001000","111111111111101101","000000000000011100","000000000000110010","111111111111001001","111111111111110011","111111111111110000","111111111111110000","111111111111100101","000000000000000111","000000000000011100","000000000000001001","111111111111111010","111111111111001011","000000000000011010","111111111111110011","111111111111111100","111111111111101010","111111111111110100","111111111111111001","111111111111111001","111111111111111001","000000000000100111","000000000000000110","000000000000100100","000000000000010100","111111111111111000","000000000000101010","111111111111011110","000000000000000001","000000000000101000","111111111111110110","000000000000011010","000000000000000000","000000000000011001","111111111111110110","000000000000010010","000000000000011001","111111111111111111","111111111111111101","000000000000000111","111111111111010100","111111111111010001","111111111111100011","000000000000000011","000000000000000111","000000000000001101"),
("111111111111101010","111111111111110000","111111111111010101","000000000000001100","111111111111111011","000000000000000000","000000000000000000","111111111111101000","000000000000011110","111111111111011100","000000000000010101","111111111111111100","000000000000010101","111111111111011001","111111111111011110","000000000000001001","111111111111101010","000000000000100001","000000000000000000","000000000000010000","111111111111101000","000000000000101110","000000000000000101","111111111111111100","111111111111111110","000000000000011010","000000000000000000","111111111111101101","000000000000001101","000000000000000110","000000000000000010","000000000000011010","000000000000001111","111111111111110100","111111111111111011","000000000000001110","111111111111101010","111111111111111101","000000000000001100","111111111111101100","000000000000100110","111111111111111110","111111111111011101","111111111111011011","000000000000011010","000000000000000101","111111111111100111","000000000000000111","111111111111111010","111111111111111011","000000000000001100","000000000000000000","000000000000011110","111111111111111100","000000000000001110","111111111111101101","111111111111110101","111111111111110111","000000000000000100","111111111111101111","000000000000011111","111111111111110100","111111111111111011","111111111111111001","111111111110111010","111111111111101000","000000000000010001","000000000000001010","111111111111110011","111111111111111110","000000000000100101","000000000000000010","000000000000000011","111111111111111110","000000000000001001","000000000000010100","111111111111111001","000000000000000001","111111111111100000","111111111111110101","111111111111111111","111111111111101100","111111111111110101","000000000000000100","000000000000100011","111111111111011100","000000000000001010","111111111111111010","111111111111101100","111111111111111100","111111111111110000","000000000000001010","111111111111110011","111111111111110101","111111111111011010","000000000000100011","000000000000011111","000000000000000101","111111111111110011","111111111111110110","000000000000000110","000000000000001010","000000000000001110","000000000000110011","111111111111110010","000000000000010101","111111111111111010","111111111111111110","000000000000100101","111111111111101100","111111111111111100","000000000000000001","000000000000000011","000000000000000111","000000000000001101","000000000000000101","111111111111110100","000000000000011011","000000000000100111","000000000000100100","111111111111101010","111111111111111110","111111111111000100","111111111111010001","111111111111101111","111111111111101011","111111111111111111","000000000000001001"),
("111111111111110011","111111111111100100","111111111111000011","000000000000001000","000000000000010111","000000000000011010","000000000000011000","111111111111100110","000000000000100011","111111111111110001","000000000000010001","000000000000000000","000000000000001001","111111111111011100","111111111111101011","000000000000010000","111111111111111100","000000000000000111","111111111111111011","000000000000001101","111111111111110011","000000000000110000","000000000000100001","111111111111110110","000000000000000001","000000000000001001","000000000000010111","111111111111111110","000000000000000111","000000000000011100","000000000000001111","000000000000011011","000000000000000000","000000000000001110","000000000000000100","000000000000000100","111111111111101001","111111111111101010","000000000000010110","000000000000001011","000000000000010000","000000000000010100","111111111111001000","111111111111101000","000000000000010010","000000000000000010","111111111111011100","000000000000001111","111111111111110100","000000000000010000","000000000000010010","000000000000001001","000000000000000110","111111111111111001","000000000000010001","000000000000000010","111111111111111111","000000000000000100","111111111111110110","000000000000001111","000000000000000110","111111111111101000","111111111111101101","000000000000000011","111111111111001101","000000000000001110","111111111111111001","000000000000100100","111111111111010001","000000000000000011","000000000000001000","000000000000010010","000000000000001001","111111111111110010","000000000000100110","000000000000010110","111111111111110110","111111111111111010","111111111111110001","000000000000000000","111111111111111101","111111111111111001","000000000000011111","111111111111110001","000000000000000110","111111111111111100","000000000000000000","000000000000010000","111111111111111000","111111111111101110","000000000000001000","111111111111110101","111111111111101100","000000000000001011","111111111111100111","000000000000001101","111111111111111001","111111111111111111","000000000000010000","000000000000010001","111111111111111100","111111111111111011","000000000000011101","000000000000001110","111111111111110010","000000000000001001","111111111111100110","000000000000001000","000000000000010110","000000000000010010","111111111111110110","000000000000101000","000000000000010010","000000000000001001","111111111111110101","000000000000100010","000000000000000110","000000000000011010","000000000000010000","000000000000011111","111111111111110001","000000000000000110","111111111111101100","111111111111010111","111111111111110010","000000000000001010","000000000000000000","111111111111111100"),
("111111111111110000","111111111111011101","111111111111011000","111111111111111101","000000000000010001","000000000000000101","000000000000011110","000000000000000101","000000000000011001","000000000000000001","000000000000100110","000000000000000111","000000000000001011","111111111111100010","111111111111001100","000000000000010010","111111111111110010","000000000000100000","000000000000000111","000000000000000000","111111111111110111","000000000000101001","000000000000000111","111111111111111101","000000000000001111","111111111111111101","111111111111111010","111111111111110100","111111111111111010","000000000000000000","111111111111110111","111111111111111000","000000000000000011","111111111111111100","000000000000010100","111111111111100011","111111111111110101","111111111111110110","111111111111111001","111111111111111100","000000000000011011","000000000000001001","111111111111011100","111111111111111010","111111111111111100","111111111111011011","000000000000000000","000000000000000100","111111111111111011","000000000000000110","000000000000001001","111111111111111101","000000000000000010","111111111111111011","000000000000000010","111111111111110111","111111111111110011","111111111111101001","000000000000000111","000000000000000111","000000000000000101","111111111111110100","000000000000000011","111111111111111100","111111111111101011","111111111111111111","000000000000001110","000000000000101100","111111111111000010","111111111111111100","111111111111111011","111111111111111001","000000000000000101","111111111111100000","000000000000100001","111111111111111111","000000000000000110","111111111111111111","000000000000010100","000000000000001011","000000000000000100","111111111111111101","111111111111110011","111111111111110010","000000000000001000","000000000000000000","000000000000000111","000000000000000011","111111111111101011","000000000000001101","000000000000000111","000000000000000101","111111111111101110","111111111111111100","000000000000001111","111111111111111000","111111111111101110","111111111111111111","111111111111111111","000000000000010100","000000000000000001","000000000000001100","000000000000010100","000000000000000101","111111111111111011","000000000000001000","111111111111100000","111111111111101000","000000000000100001","000000000000010001","111111111111101100","000000000000010101","000000000000001100","111111111111101000","111111111111110010","111111111111111011","000000000000010001","000000000000001000","000000000000000001","000000000000000100","111111111111111000","000000000000100010","000000000000010000","111111111111101101","111111111111110110","000000000000000111","000000000000000010","111111111111100110"),
("000000000000001011","111111111111111111","111111111111100001","000000000000001001","000000000000000111","000000000000000000","000000000000010100","111111111111110000","000000000000011100","000000000000000110","000000000000010001","111111111111101111","000000000000001001","000000000000000101","111111111111010110","000000000000100011","000000000000000010","000000000000010001","111111111111110101","000000000000000001","111111111111010000","111111111111111110","000000000000100010","000000000000010011","111111111111110000","000000000000001000","000000000000010000","111111111111111001","111111111111101111","000000000000001011","111111111111111011","111111111111111100","111111111111101111","000000000000001101","000000000000000000","111111111111101111","000000000000000111","000000000000001011","111111111111101101","000000000000000110","000000000000010111","000000000000001011","111111111111010110","000000000000011111","111111111111101110","111111111111110010","000000000000000001","000000000000011010","111111111111110101","000000000000000110","000000000000010000","111111111111111011","000000000000000111","000000000000000011","000000000000001001","111111111111101010","111111111111100111","000000000000001100","000000000000001101","111111111111111000","000000000000001010","000000000000000001","000000000000010100","111111111111111000","000000000000001110","000000000000011011","000000000000010101","000000000000011101","111111111111101110","000000000000100011","000000000000001001","111111111111110000","000000000000001010","111111111111110111","000000000000010100","000000000000010100","111111111111111010","111111111111111000","111111111111111000","000000000000000011","000000000000001010","111111111111100100","000000000000000100","000000000000001010","111111111111110011","111111111111011111","000000000000001101","000000000000000110","111111111111111000","111111111111110011","111111111111100011","000000000000000000","111111111111110100","000000000000011001","000000000000010010","000000000000001001","111111111111111100","111111111111110000","000000000000000001","000000000000001110","111111111111111000","111111111111111110","000000000000010010","000000000000001101","000000000000011010","000000000000000010","111111111111111010","111111111111110111","111111111111111100","000000000000001011","111111111111110001","000000000000100011","000000000000001100","111111111111101001","111111111111011100","000000000000100010","000000000000010110","000000000000011100","111111111111101101","111111111111111110","000000000000100010","000000000000001111","111111111111111100","000000000000010010","111111111111110111","000000000000000101","000000000000000010","111111111111110010"),
("111111111111111100","000000000000011000","111111111111110001","111111111111100011","000000000000010101","000000000000001000","000000000000010000","000000000000011101","111111111111111011","000000000000010101","000000000000001001","111111111111100101","111111111111111001","111111111111101010","111111111111100110","000000000000010010","000000000000000000","000000000000010010","000000000000001011","000000000000010011","111111111111100001","111111111111001111","000000000000011011","000000000000011110","111111111111110100","000000000000000010","000000000000000000","111111111111100111","111111111111110000","000000000000001111","000000000000001000","111111111111110000","111111111111111100","000000000000001000","000000000000001101","111111111111101011","000000000000010010","000000000000001001","111111111111110111","000000000000000111","000000000000100010","000000000000001111","111111111111110001","000000000000011000","000000000000010110","111111111111011111","000000000000000010","111111111111101111","000000000000001100","000000000000001010","000000000000000010","111111111111111001","000000000000001011","111111111111110110","000000000000011110","111111111111111110","111111111111100101","000000000000001001","111111111111111100","111111111111111110","111111111111111111","000000000000001110","000000000000001000","111111111111101100","111111111111111011","000000000000001101","000000000000100101","000000000000011010","111111111111010010","000000000000011101","111111111111111010","000000000000010001","000000000000001010","111111111111110000","111111111111110111","000000000000011110","000000000000010011","000000000000000111","000000000000001101","111111111111111100","000000000000001101","111111111111110111","111111111111011001","000000000000000000","000000000000010001","111111111111110000","111111111111111100","000000000000011101","111111111111111100","111111111111111111","111111111111100011","000000000000001001","000000000000010010","000000000000100101","000000000000001110","000000000000000000","111111111111111000","111111111111101110","000000000000000001","000000000000001000","111111111111111101","000000000000100100","000000000000001010","111111111111111000","000000000000000101","000000000000001010","111111111111100001","000000000000000101","000000000000001010","111111111111111010","000000000000000001","000000000000010111","000000000000010001","111111111111111001","000000000000001101","111111111111111001","000000000000010100","000000000000100111","111111111111101101","000000000000100001","000000000000010001","000000000000011100","000000000000010101","000000000000011100","111111111111011001","000000000000000011","000000000000100111","111111111111100111"),
("000000000000001010","000000000000000010","111111111111100101","000000000000000001","111111111111110110","111111111111111010","000000000000000010","111111111111110010","111111111111101000","111111111111111101","000000000000100010","111111111111101110","111111111111101100","111111111111101111","000000000000000011","000000000000011001","000000000000001100","000000000000001111","000000000000001100","000000000000010010","000000000000000011","111111111110101000","000000000000010001","111111111111111111","000000000000010001","000000000000001000","000000000000000000","000000000000001111","111111111111110011","000000000000001100","111111111111110110","111111111111110101","000000000000001001","000000000000010010","000000000000011101","000000000000000000","000000000000010101","000000000000000001","111111111111100111","111111111111110111","000000000000010001","000000000000010101","000000000000001010","000000000000010101","000000000000001011","000000000000000101","111111111111111001","000000000000010011","000000000000000001","111111111111111100","000000000000000001","111111111111110001","111111111111111001","000000000000000101","000000000000011100","111111111111101010","111111111111100011","111111111111110001","111111111111111000","111111111111111010","000000000000100101","111111111111111101","111111111111110110","000000000000000010","000000000000000111","000000000000100001","000000000000000111","000000000000100011","111111111111100110","000000000000001010","111111111111110011","000000000000010000","000000000000100010","000000000000001010","000000000000010100","000000000000011000","111111111111111111","000000000000010010","000000000000000100","000000000000010100","111111111111110111","000000000000000011","111111111111001101","000000000000000001","111111111111111010","000000000000001101","000000000000000001","000000000000000111","000000000000001100","111111111111110000","111111111111111010","000000000000001011","000000000000000000","000000000000001010","111111111111100000","111111111111111010","111111111111111010","111111111111101100","000000000000011011","000000000000010010","111111111111111100","000000000000011111","000000000000011000","111111111111101010","111111111111111101","000000000000001011","111111111111101001","000000000000001011","111111111111110011","000000000000010111","111111111111101001","000000000000100111","000000000000011011","111111111111111011","000000000000000011","000000000000000010","111111111111111001","000000000000011111","111111111111101011","000000000000001010","000000000000100100","000000000000001010","000000000000010000","000000000000011000","111111111111110011","000000000000001111","000000000000100000","111111111111100000"),
("000000000000000000","111111111111111110","111111111111101101","111111111111110001","000000000000001000","111111111111111100","111111111111111100","111111111111110111","111111111111111100","000000000000001001","000000000000010011","000000000000000101","111111111111110011","111111111111010010","000000000000010000","000000000000110010","111111111111111001","000000000000011000","111111111111110110","000000000000001111","111111111111101110","111111111110100100","111111111111110101","111111111111110010","111111111111111101","000000000000000100","111111111111110110","000000000000010000","111111111111111110","000000000000000010","111111111111111011","000000000000001000","000000000000000001","000000000000001010","000000000000011011","000000000000001001","000000000000000000","111111111111111100","111111111111010011","111111111111111111","000000000000100011","111111111111110110","000000000000000110","000000000000001011","111111111111111001","111111111111111010","000000000000011101","000000000000101001","000000000000000100","111111111111110111","000000000000000100","000000000000001011","111111111111111110","111111111111111000","000000000000000000","111111111111110011","111111111111100101","000000000000000000","000000000000000100","000000000000000100","000000000000010101","000000000000000000","000000000000000011","000000000000000110","111111111111111110","111111111111111011","000000000000001100","000000000000100111","111111111111101010","111111111111101100","000000000000000000","000000000000001011","111111111111111110","000000000000001101","111111111111110111","000000000000011011","111111111111110000","000000000000000000","000000000000000000","111111111111111010","000000000000000000","000000000000000111","111111111111011101","111111111111110101","111111111111111100","000000000000000000","000000000000011001","000000000000001101","000000000000010010","111111111111100101","111111111111111000","000000000000000001","000000000000001001","000000000000000111","111111111111111101","000000000000000000","000000000000000000","111111111111110110","000000000000001111","000000000000000101","111111111111110100","000000000000010001","000000000000011111","000000000000011010","111111111111101111","111111111111111011","111111111111101101","000000000000000110","111111111111100000","000000000000011100","111111111111100000","000000000000011101","000000000000011100","111111111111111101","111111111111111111","000000000000010010","000000000000000111","000000000000110000","111111111111111011","000000000000011001","000000000000100101","111111111111111101","000000000000010110","000000000000010111","111111111111011010","000000000000010110","000000000000001100","111111111111111110"),
("000000000000010100","111111111111110101","000000000000001000","111111111111111010","000000000000000001","000000000000011010","111111111111100010","111111111111110111","111111111111111011","000000000000000011","000000000000011101","111111111111101100","111111111111101101","111111111111100110","000000000000011010","000000000000100011","111111111111111110","000000000000000000","000000000000010001","000000000000000010","111111111111101010","111111111111000101","000000000000010010","111111111111101000","111111111111101101","000000000000011001","111111111111100100","000000000000000010","000000000000000000","000000000000010101","111111111111100001","000000000000001010","000000000000000010","000000000000010011","000000000000001111","111111111111110111","111111111111101101","000000000000001000","111111111111011110","000000000000001101","000000000000011001","000000000000001001","000000000000101100","111111111111111101","000000000000001010","000000000000010010","000000000000000001","000000000000100100","111111111111111010","111111111111110101","111111111111101101","111111111111100000","000000000000000010","111111111111111011","000000000000000100","111111111111111111","111111111111110010","000000000000001001","000000000000001001","111111111111101101","000000000000001100","000000000000001000","111111111111100101","111111111111101110","111111111111100010","111111111111101000","000000000000100011","000000000000101001","111111111111101010","000000000000000110","000000000000011110","111111111111111001","111111111111111100","000000000000000000","000000000000011010","111111111111110110","000000000000001000","111111111111111111","111111111111111000","111111111111111110","111111111111111110","000000000000000101","111111111111011100","111111111111111100","000000000000101100","111111111111111100","111111111111110101","000000000000000101","111111111111110011","111111111111101100","000000000000010101","000000000000000100","000000000000100010","000000000000001110","111111111111101101","000000000000001011","000000000000000110","111111111111110100","000000000000110000","111111111111101100","000000000000010111","000000000000011000","000000000000001100","000000000000000010","111111111111100011","000000000000001001","000000000000001000","000000000000100011","111111111111100111","111111111111101110","111111111111110111","000000000000010110","000000000000010011","000000000000001100","000000000000000000","000000000000011110","000000000000001001","000000000000001001","111111111111101010","000000000000010010","000000000000100011","111111111111100000","111111111111110110","000000000000110010","111111111111000011","000000000000010001","000000000000011100","000000000000000110"),
("111111111111111111","000000000000000000","000000000000000111","111111111111111011","111111111111111100","000000000000010010","111111111111100011","000000000000010011","111111111111110001","000000000000000100","000000000000011110","000000000000010101","111111111111110110","111111111111011011","000000000000010101","000000000000010111","000000000000000000","000000000000011001","111111111111111010","111111111111111110","111111111111110000","111111111111100011","000000000000000101","111111111111100010","111111111111110100","111111111111110100","111111111111101001","111111111111110110","000000000000001111","000000000000100110","111111111111101001","000000000000101010","111111111111101110","000000000000001101","000000000000001001","000000000000010110","111111111111110000","000000000000001111","111111111111110110","111111111111110011","000000000000101011","111111111111111101","000000000000010111","000000000000000010","111111111111111011","000000000000011010","111111111111110111","000000000000000101","000000000000010110","000000000000000000","111111111111101001","000000000000001110","111111111111110111","111111111111110010","000000000000001001","111111111111101110","000000000000011001","000000000000001110","000000000000000111","000000000000000000","000000000000010000","000000000000001000","111111111111101011","111111111111111110","111111111111111000","000000000000001001","000000000000000001","000000000000110001","111111111111111100","000000000000000100","000000000000001110","111111111111111000","111111111111111110","000000000000001101","000000000000000010","111111111111100011","111111111111110000","111111111111111110","000000000000000011","000000000000000010","111111111111111110","000000000000000101","111111111111101100","111111111111110011","000000000000011000","111111111111100011","000000000000100010","000000000000010101","111111111111111110","000000000000000011","000000000000100101","111111111111111111","000000000000000010","111111111111111000","000000000000000001","000000000000001101","000000000000001000","000000000000001010","000000000000001101","111111111111100010","000000000000001001","000000000000001001","000000000000010011","000000000000011111","111111111111111111","111111111111110111","000000000000001100","000000000000000101","111111111111101111","111111111111100111","000000000000000010","000000000000101011","000000000000100101","111111111111111110","111111111111111100","111111111111110111","000000000000000100","000000000000001010","111111111111111111","000000000000010111","000000000000010101","000000000000000100","111111111111111011","000000000000011111","111111111111101111","000000000000011000","000000000000010110","111111111111111000"),
("111111111111111101","000000000000000010","000000000000000101","000000000000010011","000000000000001011","000000000000000000","111111111111011100","111111111111101101","111111111111101111","000000000000000010","000000000000010111","000000000000010010","000000000000010110","111111111111010110","000000000000010101","000000000000100001","111111111111110100","111111111111111111","111111111111100100","000000000000000110","000000000000000011","000000000000001111","000000000000000110","111111111111101100","111111111111101100","000000000000001111","111111111111110000","000000000000001111","000000000000001000","000000000000000101","000000000000001101","000000000000000110","111111111111110000","000000000000010010","111111111111111101","000000000000011110","000000000000001110","000000000000010001","000000000000000010","000000000000000000","000000000000011001","111111111111100011","000000000000000101","111111111111110101","000000000000000011","000000000000000000","000000000000000000","111111111111101111","111111111111110100","000000000000000111","111111111111101001","000000000000000000","111111111111101111","000000000000000000","111111111111101100","111111111111110001","000000000000010100","000000000000010010","111111111111111011","111111111111111101","111111111111111111","000000000000010001","111111111111111100","111111111111101000","111111111111110011","111111111111111011","111111111111011111","000000000000001111","000000000000000000","000000000000000001","000000000000010101","000000000000001110","111111111111101110","000000000000000110","000000000000001010","111111111111011001","111111111111110111","000000000000000100","111111111111110011","111111111111101101","000000000000010011","000000000000010101","111111111111100001","111111111111100101","111111111111111011","000000000000000101","000000000000011010","000000000000001111","000000000000010111","000000000000010000","000000000000011110","000000000000001010","000000000000000000","111111111111100100","000000000000010111","111111111111101110","000000000000010001","111111111111110000","000000000000010101","111111111111010100","000000000000000011","000000000000001101","000000000000011111","000000000000000000","111111111111101001","111111111111111101","111111111111110010","000000000000000101","000000000000001111","111111111111100001","111111111111111110","000000000000110101","000000000000010110","000000000000001010","000000000000000110","000000000000000100","111111111111110111","000000000000000101","000000000000010001","000000000000010000","111111111111111111","000000000000010011","111111111111110111","000000000000010111","111111111111100100","111111111111111100","111111111111110111","000000000000001111"),
("000000000000100101","000000000000001010","111111111111100111","000000000000000101","000000000000011011","000000000000010001","111111111111110100","111111111111100010","111111111111110110","111111111111111011","000000000000001101","000000000000100000","000000000000010100","111111111111100000","000000000000001100","000000000000000111","000000000000010100","111111111111110111","111111111111110100","111111111111110111","000000000000000111","000000000000010101","000000000000001100","111111111111110111","111111111111100110","000000000000001001","000000000000000101","000000000000011000","000000000000000011","000000000000010100","111111111111111110","111111111111111100","000000000000000100","000000000000000000","111111111111110111","000000000000011111","111111111111101100","000000000000010110","000000000000000111","000000000000000101","000000000000001010","111111111111101101","111111111111100011","111111111111111111","000000000000011101","111111111111101100","000000000000010010","000000000000010011","111111111111111110","000000000000001010","111111111111111000","000000000000010000","111111111111101010","111111111111111101","111111111111111111","111111111111111111","000000000000011100","000000000000000110","000000000000000000","111111111111101100","000000000000001100","000000000000010001","111111111111101000","111111111111101111","111111111111001111","111111111111101101","111111111111101000","000000000000010111","111111111111110111","111111111111111110","000000000000000011","000000000000010100","111111111111110001","111111111111101110","000000000000011110","111111111111011100","111111111111111110","000000000000001110","000000000000000110","111111111111011011","000000000000001010","000000000000010011","111111111111110010","111111111111011111","000000000000100000","111111111111010001","000000000000001001","000000000000000110","000000000000100000","111111111111110111","000000000000010110","111111111111111000","000000000000010101","111111111111101010","000000000000010101","111111111111110000","000000000000001101","000000000000001010","000000000000000010","111111111111101100","000000000000011111","000000000000001010","000000000000010000","000000000000010101","111111111111111010","111111111111110010","111111111111110010","111111111111101111","000000000000000111","111111111111011110","111111111111110111","000000000000101100","000000000000010100","000000000000000110","000000000000000001","000000000000010001","111111111111110110","000000000000000010","000000000000000110","000000000000001000","000000000000001011","111111111111110100","111111111111101111","000000000000101101","111111111111100110","000000000000000011","000000000000000101","000000000000001011"),
("000000000000010101","000000000000100100","111111111111101000","000000000000010110","111111111111111011","000000000000011000","111111111111101001","000000000000000111","111111111111110110","000000000000001101","000000000000101001","000000000000001011","000000000000010000","111111111111011110","000000000000000000","000000000000100001","000000000000010001","111111111111111111","111111111111111100","000000000000010000","111111111111011101","000000000000010011","111111111111111110","111111111111011110","111111111111111001","000000000000000111","000000000000000011","000000000000000000","000000000000000100","111111111111110111","000000000000010000","000000000000001111","111111111111111100","000000000000011111","111111111111110101","000000000000010000","111111111111101111","000000000000011000","000000000000000100","000000000000001010","000000000000010110","111111111111110010","000000000000000000","111111111111111111","000000000000000000","111111111111110111","111111111111110110","000000000000011011","111111111111101100","111111111111101100","111111111111101000","111111111111101011","111111111111110110","000000000000000110","111111111111110100","111111111111110111","111111111111111101","111111111111110010","111111111111111000","111111111111110101","111111111111111111","111111111111111111","000000000000000111","111111111111110000","111111111111101010","111111111111110000","111111111110111000","000000000000100101","111111111111110110","111111111111110111","000000000000100110","000000000000000011","000000000000000011","111111111111101100","000000000000011000","111111111111110000","000000000000010101","000000000000010000","111111111111110011","111111111111100100","111111111111110100","000000000000001001","111111111111110100","111111111110110001","000000000000011010","111111111111101011","111111111111110110","000000000000000000","000000000000001010","000000000000011000","000000000000001101","111111111111110110","111111111111101100","000000000000000010","111111111111100111","111111111111001110","111111111111101110","000000000000001011","111111111111110101","111111111111111111","000000000000000010","000000000000010011","111111111111101011","000000000000010011","111111111111100011","111111111111110110","111111111111101001","111111111111111100","000000000000001110","111111111111101010","111111111111111110","000000000000100111","000000000000100000","111111111111100101","111111111111101001","000000000000011000","000000000000001001","000000000000001000","111111111111111011","000000000000100100","000000000000100000","000000000000000000","111111111111111011","000000000000111001","111111111111111100","111111111111111001","000000000000000001","000000000000010111"),
("000000000000101001","000000000000100010","111111111111101110","000000000000011110","000000000000001000","000000000000101001","111111111111011111","111111111111111011","111111111111101110","000000000000001100","000000000000111001","000000000000010000","000000000000000111","111111111111101001","000000000000000000","000000000000000010","000000000000100001","000000000000100100","000000000000000001","000000000000011011","111111111111111100","000000000000001001","000000000000001111","111111111111101101","111111111111100110","000000000000011001","111111111111111010","111111111111111111","000000000000000111","111111111111110011","000000000000001010","000000000000001011","111111111111110000","111111111111111010","000000000000000100","000000000000011100","111111111111011101","111111111111111110","111111111111110000","000000000000010110","000000000000010011","000000000000001000","111111111111111000","000000000000000011","000000000000011100","111111111111110111","111111111111110110","000000000000000000","000000000000001011","111111111111101111","111111111111100001","111111111111111101","111111111111100111","000000000000011011","000000000000000000","111111111111101111","111111111111100111","111111111111111110","111111111111011111","111111111111110000","111111111111101000","000000000000010011","111111111111110110","111111111111111000","111111111111100001","111111111111011011","111111111110001011","000000000000010110","111111111111110101","000000000000001100","000000000000010100","000000000000000110","111111111111011010","111111111111110011","000000000000101101","111111111111100011","000000000000000100","000000000000100001","111111111111100001","000000000000000100","111111111111110100","000000000000000001","111111111111111101","111111111110110000","000000000000001100","111111111111010011","111111111111111011","000000000000010000","111111111111110001","000000000000010101","000000000000000110","111111111111111010","111111111111100101","000000000000000000","000000000000000110","111111111111001110","000000000000001010","000000000000001000","111111111111011011","111111111111110110","000000000000000001","000000000000000111","111111111111011010","111111111111111111","111111111111100111","000000000000000100","111111111111101101","111111111111101101","000000000000000000","111111111111011111","111111111111110100","000000000000101000","000000000000011101","111111111111111110","000000000000000011","000000000000000000","111111111111111101","111111111111110001","111111111111001011","000000000000010000","000000000000000100","111111111111111010","000000000000001111","000000000000011100","111111111111010101","111111111111110100","000000000000001001","111111111111101110"),
("000000000000101010","000000000000101110","111111111111101010","000000000000000011","000000000000011100","000000000000010111","111111111111010001","000000000000001000","000000000000001100","111111111111111011","000000000000010111","000000000000110000","000000000000001110","000000000000001001","111111111111100101","000000000000000011","000000000000010111","000000000000000110","111111111111101101","111111111111111001","000000000000001101","111111111111011010","000000000000010111","111111111111110011","111111111111101011","000000000000000000","000000000000001000","111111111111111001","111111111111110010","111111111111111010","000000000000001101","111111111111110110","111111111111110100","000000000000000000","111111111111110111","000000000000010010","111111111111011111","111111111111111101","000000000000000100","000000000000001010","000000000000011010","111111111111111010","000000000000000100","000000000000001011","000000000000010100","111111111111010110","111111111111100110","000000000000001100","111111111111111110","111111111111100011","000000000000001000","000000000000000110","000000000000000100","000000000000100110","000000000000001000","000000000000001101","111111111111100111","111111111111011001","111111111111100101","111111111111110011","111111111111001011","000000000000100001","000000000000001010","111111111111101000","111111111111110100","000000000000000000","111111111110101100","000000000000001101","000000000000000101","111111111111110000","000000000000010001","000000000000001001","111111111110101001","111111111111101110","000000000000101110","111111111111100100","111111111111110010","111111111111111010","111111111111100110","111111111111110110","111111111111101101","111111111111111000","111111111111111101","111111111111011011","000000000000010001","111111111111011000","000000000000001000","111111111111111011","000000000000000000","111111111111110110","111111111111111100","111111111111110001","000000000000000110","000000000000000100","111111111111110001","111111111111000001","111111111111101010","111111111111110000","111111111111110000","000000000000000111","000000000000000000","000000000000010110","111111111111100000","000000000000101001","111111111111110001","111111111111100111","111111111111110000","111111111111101001","000000000000001001","111111111111100000","000000000000000011","000000000000010001","000000000000001010","000000000000000001","000000000000000111","111111111111011110","111111111111011111","111111111111101101","111111111111010011","000000000000000000","000000000000001001","111111111111111010","111111111111101101","000000000000001010","111111111111011001","000000000000010110","111111111111111011","000000000000001010"),
("000000000000100010","000000000000001001","000000000000000100","111111111111111111","000000000000011101","000000000000001010","000000000000000101","000000000000100111","111111111111111000","111111111111111100","000000000000000111","000000000000011100","000000000000010110","000000000000100001","111111111111100101","000000000000011011","000000000000010010","000000000000000011","111111111111100100","000000000000000100","000000000000000000","111111111111110011","111111111111111100","111111111111011101","111111111111010110","000000000000001100","111111111111111111","111111111111111011","000000000000001011","111111111111100101","000000000000010000","111111111111101000","111111111111100010","000000000000010101","000000000000010100","111111111111110010","000000000000000000","000000000000011001","111111111111111000","111111111111101011","000000000000100001","000000000000000000","111111111111101001","111111111111110111","000000000000010100","111111111111010110","111111111111000000","000000000000010000","000000000000001010","111111111111110111","000000000000000100","000000000000010101","111111111111011010","000000000000100001","000000000000001011","000000000000000101","111111111111101001","111111111111001111","111111111111111000","111111111111111000","111111111111000001","000000000000010011","111111111111111101","111111111111110110","000000000000010011","111111111111100001","111111111110110101","111111111111011000","111111111111110011","111111111111101100","000000000000000011","111111111111110001","111111111110101110","111111111111101111","000000000000001011","111111111111111100","000000000000001010","000000000000000000","111111111111110000","111111111111111001","111111111111100100","111111111111111001","000000000000010011","111111111111100000","000000000000001111","111111111111111001","111111111111111011","000000000000001110","111111111111101110","111111111111101101","111111111111110010","111111111111010110","111111111111111110","111111111111111111","111111111111011111","111111111111010110","111111111111100011","111111111111110100","111111111110111001","111111111111111011","000000000000001001","111111111111111101","111111111111010110","000000000000000000","111111111111101110","111111111111111101","111111111111111001","111111111111000010","111111111111111101","111111111111011011","111111111111111000","000000000000000000","111111111111110101","000000000000000110","000000000000001000","111111111111101000","111111111111010111","000000000000010101","111111111111101110","000000000000000010","000000000000000011","111111111111110010","111111111111111010","111111111111111100","111111111111100000","111111111111111001","000000000000000101","000000000000001011"),
("000000000000010010","000000000000001011","000000000000001101","000000000000001010","000000000000001101","000000000000001111","000000000000000000","000000000000100101","000000000000001000","000000000000001011","000000000000011010","000000000000000110","000000000000011010","000000000000000001","111111111111011110","000000000000001001","111111111111110101","000000000000001010","111111111111111101","000000000000100011","111111111111110011","111111111111100001","111111111111111110","111111111111110011","111111111111100011","000000000000000101","000000000000011010","000000000000011010","000000000000000100","111111111111111001","000000000000011101","111111111111011110","000000000000000000","111111111111110111","000000000000000011","000000000000000010","000000000000000101","000000000000100010","111111111111100100","111111111111100110","000000000000000001","111111111111110011","111111111111110010","111111111111111011","000000000000101001","111111111111100111","111111111111001010","000000000000011000","000000000000000111","111111111111110000","111111111111110001","000000000000001100","111111111111110001","111111111111111000","111111111111101000","000000000000000110","111111111111011101","111111111111011110","111111111111100010","111111111111111010","111111111110111100","000000000000000000","000000000000011010","000000000000000111","000000000000000001","000000000000001000","111111111111101100","000000000000000111","111111111111101111","000000000000000101","000000000000000101","000000000000000000","111111111111010011","111111111111110110","000000000000001110","111111111111111001","000000000000010001","111111111111100111","111111111111111000","000000000000000011","111111111111100100","000000000000010101","000000000000011011","111111111111100101","000000000000001111","111111111111101100","000000000000000101","000000000000001110","000000000000011101","111111111111110011","000000000000001111","111111111111111101","000000000000001100","111111111111101100","111111111111100101","111111111111101011","111111111111110011","000000000000001001","111111111111010010","111111111111111100","000000000000010111","000000000000010000","111111111110101110","000000000000000111","111111111111100100","111111111111111001","000000000000001010","111111111111011110","111111111111100010","111111111111101100","111111111111110010","000000000000001100","000000000000100011","000000000000000100","000000000000100110","000000000000000010","111111111111110011","000000000000011101","111111111111011111","000000000000001001","000000000000010100","111111111111110111","111111111111101000","000000000000000001","111111111111010010","000000000000000001","000000000000000000","111111111111101001"),
("000000000000110001","111111111111101000","111111111111111110","000000000000011111","111111111111111000","000000000000001101","000000000000010000","000000000000111101","000000000000001100","111111111111110011","000000000000001101","000000000000001001","000000000000101011","111111111111111111","111111111111110101","000000000000100101","000000000000001010","000000000000011100","111111111111110011","000000000000011010","111111111111111011","111111111111000100","111111111111110101","111111111111100111","111111111111111000","000000000000010010","000000000000100001","000000000000000010","000000000000000101","111111111111100101","000000000000110100","111111111111011001","111111111111101101","000000000000001010","111111111111110001","111111111111010111","111111111111111110","000000000000001111","111111111111110101","111111111111011111","000000000000100100","111111111111101101","000000000000000001","000000000000001110","000000000000010100","111111111111110100","111111111110111011","000000000000010100","111111111111111011","111111111111011100","111111111111111100","000000000000000011","111111111111011101","000000000000010001","111111111111111101","000000000000100010","111111111111011101","111111111111011011","111111111111011100","111111111111111100","111111111111011010","000000000000000011","111111111111111110","111111111111110001","000000000000011010","000000000000000010","111111111111110000","111111111111101000","111111111111100010","111111111111100101","111111111111111111","111111111111110100","111111111111101110","111111111111100100","111111111111100010","000000000000001100","000000000000100110","000000000000001100","111111111111110000","000000000000001101","111111111111111111","000000000000000010","000000000000000101","111111111111011111","111111111111111100","111111111111111110","000000000000010110","000000000000000010","000000000000010110","111111111111001011","111111111111111011","111111111111101110","111111111111110110","111111111111100110","111111111111111011","000000000000001101","000000000000011110","111111111111111010","111111111111010011","111111111111101110","000000000000100111","111111111111110001","111111111111100000","000000000000011011","000000000000000000","111111111111101101","111111111111101100","111111111111010111","111111111111110001","111111111111100010","111111111111111001","000000000000011001","111111111111111111","111111111111010011","111111111111111110","111111111111100011","111111111111001111","000000000000100000","111111111111100111","111111111111110010","000000000000010110","111111111111110110","111111111111101110","000000000000010001","111111111111110010","000000000000000101","111111111111111110","111111111111101001"),
("000000000000011000","000000000000011010","000000000000010000","000000000000011010","000000000000010001","111111111111111101","000000000000001110","111111111111100110","111111111111011110","111111111111100011","000000000000100110","111111111111101011","000000000001001000","000000000000100110","000000000000000101","000000000000001110","111111111111110011","000000000000000111","111111111111001011","111111111111101111","000000000000011100","111111111111110111","000000000000001101","111111111111111000","111111111111110101","000000000000001100","000000000000000111","000000000000010110","000000000000000110","111111111111011011","000000000000111000","111111111111101100","111111111111101111","000000000000000110","000000000000100000","111111111111110101","111111111111111011","000000000000011110","111111111111101111","000000000000000001","000000000000000111","111111111111101011","111111111111110101","000000000000001000","111111111111110010","000000000000010000","111111111111010000","111111111111101010","111111111111101110","111111111111001111","111111111111011111","111111111111101101","111111111111101101","000000000001000001","000000000000100111","000000000000001110","111111111111101111","111111111111101110","111111111111110100","000000000000001100","111111111111001111","000000000000110010","000000000000000111","111111111111100111","000000000000101010","111111111111110001","111111111111101010","111111111111011000","000000000000001011","111111111111110100","111111111111110110","000000000000001110","111111111111110110","111111111111110100","111111111111111100","111111111111111011","000000000000001001","111111111111110111","000000000000010011","111111111111101101","000000000000010010","000000000000000000","000000000000001100","111111111111110110","000000000000011100","111111111111111111","000000000000011111","111111111111111100","111111111111100111","111111111111101000","111111111111111011","111111111111101000","111111111111101001","111111111111110111","000000000000011010","111111111111110010","000000000000000010","000000000000010000","000000000000011001","111111111111100101","111111111111111001","111111111111100100","111111111111100101","111111111111111000","111111111111111100","111111111111110111","000000000000001110","111111111111110010","111111111111011010","111111111111110001","000000000000000100","000000000000110111","111111111110111100","111111111111100000","000000000000001110","111111111111100011","111111111111000011","000000000000000110","000000000000000000","111111111111101110","000000000000010001","000000000000010100","000000000000100110","000000000000100011","000000000000010010","111111111111111101","000000000000010000","111111111111110011"),
("000000000000100101","111111111111111111","000000000000100010","111111111111111111","000000000000001100","111111111111111000","111111111111110111","000000000000000000","000000000000001110","111111111111001111","000000000000010110","111111111111111100","000000000000010111","000000000000100001","111111111111101110","000000000000001011","111111111111110001","000000000000001110","111111111111111011","000000000000010010","000000000000111010","111111111111111010","111111111111110011","111111111111111111","000000000000000000","000000000000001001","111111111111101111","111111111111111011","000000000000010100","111111111111101001","000000000000100101","000000000000001011","111111111111110101","000000000000010010","000000000000011010","000000000000000000","000000000000001110","000000000000100110","111111111111100010","111111111111101100","111111111111110101","111111111111010101","111111111111111101","111111111111110011","111111111111111010","111111111111110011","111111111111101110","000000000000011111","111111111111110101","111111111111101100","111111111111110000","000000000000001101","111111111111110010","000000000000101000","000000000000011011","111111111111111011","111111111111111110","111111111111101110","111111111111010010","111111111111111111","111111111111101000","000000000000000011","000000000000000011","111111111111011100","000000000000000100","000000000000001100","000000000000001001","000000000000000000","000000000000101101","000000000000000010","111111111111111011","111111111111111111","111111111111111110","111111111111111000","000000000000000000","111111111111110110","111111111111110111","000000000000100000","111111111111110100","111111111111110111","000000000000000100","000000000000000111","111111111111110000","111111111111001110","000000000000001101","000000000000001110","111111111111110110","000000000000001101","111111111111010001","000000000000010100","000000000000010110","111111111111101100","000000000000011000","111111111111110101","111111111111011110","000000000000010010","111111111111101110","111111111111011111","111111111111101111","000000000000000000","000000000000000110","000000000000001100","111111111111110010","000000000000000101","111111111111110001","111111111111011101","000000000000000110","111111111111101010","000000000000001011","111111111111011111","000000000000000000","000000000000010100","111111111111101100","111111111111000111","111111111111101011","111111111111101011","111111111111110001","111111111111111101","111111111111111110","111111111111111011","000000000000011001","000000000000100000","111111111111110101","000000000000010110","111111111111110001","000000000000100001","000000000000100000","111111111111110000"),
("111111111111101011","000000000000001011","111111111111011100","000000000000001100","000000000000101011","111111111111011101","000000000000001000","111111111111110111","111111111111110001","000000000000011011","000000000000011111","111111111111111100","111111111111101111","111111111111100111","111111111111110000","000000000000100100","000000000000101001","000000000000001110","111111111111010110","000000000000010101","111111111111010111","111111111111101101","000000000000011111","000000000000000010","000000000000011001","111111111111011001","111111111111110111","111111111111111100","000000000000001101","111111111111110110","111111111111100100","111111111111011101","000000000000100001","000000000000001000","000000000000001110","000000000000000110","000000000000011101","000000000000100001","111111111111110001","111111111111111101","111111111111101101","111111111111101110","000000000000001011","000000000000101100","111111111111101110","111111111111111000","000000000000001001","000000000000100001","000000000000001010","111111111111000100","000000000000000000","000000000000101111","000000000000000011","111111111111110110","111111111111101110","111111111111101100","111111111111101110","000000000000010001","000000000000001101","111111111111101101","111111111111111101","000000000000100110","000000000000010101","111111111111101110","000000000000100100","000000000000000010","000000000000100101","000000000000011110","000000000000010010","000000000000000101","111111111111101000","111111111111110010","111111111111101000","000000000000001100","111111111111100010","000000000000011011","111111111111100001","111111111111110011","111111111111100001","000000000000100100","000000000000100001","111111111111101000","000000000000001111","000000000000000000","000000000000000011","000000000000110011","000000000000010011","000000000000100001","111111111111010101","111111111111101101","000000000000011010","111111111111101111","000000000000010110","000000000000110010","111111111111000111","000000000000000001","000000000000010101","111111111111101110","000000000000001101","111111111111010110","111111111111100110","000000000000001001","000000000000001010","111111111111101011","111111111111111101","000000000000011111","111111111111110001","111111111111101010","000000000000000001","000000000000100100","111111111111000110","000000000000011000","000000000000000111","111111111111110110","111111111111011000","000000000000001011","111111111111111101","000000000000100001","111111111111110000","000000000000000000","000000000000100111","000000000000011110","111111111111101010","000000000000010111","000000000000010100","111111111111110100","000000000000000110","111111111111010100"),
("111111111111111011","000000000000001101","000000000000010010","111111111111111010","000000000000000111","111111111111110010","111111111111111111","000000000000001001","000000000000000000","111111111111111110","000000000000000011","111111111111111000","111111111111110100","000000000000000000","111111111111110101","111111111111110101","111111111111101110","111111111111110111","000000000000001000","111111111111111111","000000000000001000","000000000000001100","111111111111111011","000000000000001000","111111111111111001","000000000000001010","111111111111111000","111111111111111011","111111111111101100","111111111111101101","111111111111101111","111111111111101110","000000000000000010","000000000000000101","111111111111110101","111111111111110101","000000000000000100","111111111111111010","111111111111110100","000000000000001000","000000000000000011","000000000000000101","000000000000000011","000000000000001101","000000000000000111","111111111111111111","000000000000010001","111111111111110111","000000000000010000","000000000000000000","111111111111111001","111111111111110010","000000000000000110","111111111111111000","111111111111111100","000000000000001000","111111111111110101","000000000000000001","000000000000000000","111111111111111001","111111111111110101","000000000000001111","111111111111110101","111111111111111111","111111111111111100","000000000000001010","000000000000010100","000000000000001001","000000000000000000","000000000000000100","000000000000001101","000000000000001110","000000000000010010","111111111111110111","000000000000000000","111111111111101111","111111111111110001","111111111111110000","000000000000010000","111111111111101101","111111111111110011","111111111111101100","000000000000010000","111111111111110111","000000000000001100","111111111111111100","111111111111111110","000000000000010100","000000000000000110","111111111111110100","000000000000010011","000000000000000110","111111111111111000","000000000000000000","111111111111111001","111111111111101100","000000000000000000","111111111111110100","111111111111111110","111111111111110000","111111111111110101","111111111111111001","000000000000000111","000000000000010001","111111111111101110","111111111111110010","000000000000001110","000000000000001110","111111111111111111","111111111111111011","000000000000001110","111111111111101111","000000000000010001","000000000000001100","000000000000001011","000000000000000110","111111111111110111","111111111111101100","111111111111111100","000000000000000011","111111111111110111","111111111111111000","111111111111111110","111111111111111010","000000000000000101","111111111111111001","111111111111110110","000000000000001001"),
("000000000000000010","111111111111111000","000000000000000011","000000000000001011","000000000000001101","111111111111111011","111111111111111111","000000000000000100","111111111111111110","111111111111111110","000000000000000001","000000000000010001","111111111111110110","000000000000011010","111111111111111100","111111111111101101","000000000000010001","000000000000001011","000000000000001110","111111111111101001","111111111111110110","111111111111110101","111111111111111011","000000000000000000","000000000000001011","000000000000000000","111111111111111101","000000000000010000","111111111111111101","000000000000010001","000000000000000110","111111111111110101","111111111111100111","000000000000010111","000000000000010100","000000000000001100","111111111111110010","111111111111110010","111111111111101101","111111111111110110","111111111111110101","000000000000010011","000000000000000000","000000000000010000","111111111111111110","000000000000010011","000000000000010100","111111111111101111","000000000000000101","111111111111110110","000000000000001101","111111111111101011","111111111111110001","000000000000010010","000000000000000001","111111111111111101","000000000000001001","111111111111101011","000000000000001111","111111111111111110","111111111111101101","111111111111111101","111111111111111000","000000000000010000","111111111111110110","000000000000000111","000000000000001100","111111111111111011","111111111111111011","000000000000000110","000000000000000011","111111111111110010","000000000000001011","111111111111111101","000000000000010010","111111111111110100","111111111111110111","000000000000000101","111111111111101011","111111111111101000","111111111111110010","111111111111101101","000000000000010001","000000000000000001","000000000000010001","000000000000000000","111111111111110000","000000000000010101","111111111111111011","000000000000010011","000000000000010011","111111111111101010","000000000000000010","000000000000010101","111111111111111010","111111111111110011","111111111111110110","111111111111100110","000000000000000100","000000000000000110","111111111111111001","111111111111111110","000000000000001000","111111111111110101","111111111111111100","000000000000010001","111111111111110111","111111111111111100","111111111111101111","000000000000000000","111111111111101100","111111111111111001","000000000000000000","111111111111110011","000000000000001110","111111111111110011","000000000000001001","000000000000000001","000000000000001011","111111111111110000","111111111111110101","000000000000000110","111111111111111000","000000000000001111","000000000000001111","000000000000000111","000000000000000011","000000000000000001"),
("000000000000000010","111111111111111110","111111111111110101","111111111111111011","111111111111110100","111111111111111101","000000000000000100","000000000000010000","000000000000001001","000000000000000011","000000000000000001","111111111111101100","111111111111110000","111111111111110000","000000000000000000","000000000000000110","111111111111111011","111111111111111100","111111111111110010","000000000000010011","111111111111111100","000000000000001100","000000000000001000","111111111111101101","111111111111111001","111111111111111001","111111111111110101","000000000000001000","111111111111111011","111111111111110000","000000000000000111","111111111111110101","111111111111110100","000000000000001010","111111111111111100","000000000000010011","111111111111101111","111111111111111100","000000000000001100","000000000000001111","000000000000001110","111111111111111000","111111111111101111","000000000000010101","111111111111111101","000000000000001111","000000000000010010","000000000000000100","000000000000000110","000000000000001010","000000000000010101","000000000000000101","000000000000001100","111111111111111001","000000000000000000","111111111111101100","111111111111111100","000000000000010111","000000000000001111","000000000000000101","000000000000010101","000000000000001100","111111111111110011","000000000000000101","000000000000000000","111111111111111011","000000000000000000","000000000000000111","000000000000010111","000000000000000111","000000000000010001","000000000000010000","000000000000001000","111111111111111011","000000000000000111","000000000000010101","111111111111101100","111111111111110011","111111111111111000","000000000000000000","000000000000001001","000000000000001000","000000000000001101","000000000000010111","000000000000010010","111111111111110101","111111111111111000","000000000000010001","111111111111101111","111111111111111110","111111111111110001","000000000000000111","111111111111110101","000000000000001001","111111111111111010","000000000000001001","111111111111110111","111111111111111010","111111111111110110","111111111111110011","000000000000001001","000000000000001101","000000000000001000","000000000000000001","111111111111101100","111111111111111110","111111111111110001","000000000000000001","000000000000001110","111111111111110110","111111111111110100","000000000000001000","111111111111101110","111111111111110111","111111111111110010","000000000000010111","000000000000001110","000000000000000001","000000000000001100","111111111111110111","111111111111110001","111111111111111010","000000000000001100","000000000000010001","000000000000000000","000000000000000000","111111111111110000","111111111111111000"),
("111111111111111000","111111111111111111","111111111111011101","000000000000011010","111111111111101110","000000000000011011","000000000000000110","000000000000011111","000000000000010011","111111111111110001","000000000000001010","111111111111110010","000000000000011000","111111111111111011","111111111111101111","000000000000011110","000000000000110110","111111111111111001","111111111111111011","000000000000010011","111111111111111110","111111111111101101","000000000000001110","111111111111001110","111111111111100100","000000000000101011","000000000000001011","000000000000101100","000000000000000011","111111111111100100","111111111111111000","111111111111101111","000000000000001101","111111111111101110","111111111111101100","111111111111110010","111111111111110110","111111111111111001","111111111111111010","111111111111101010","111111111111100011","111111111111100011","000000000000000100","000000000000001001","111111111111111110","000000000000001011","111111111111110001","111111111111110001","111111111111111010","111111111111111011","000000000000000011","000000000000101001","111111111111011100","111111111111110000","000000000000010110","000000000000000101","111111111111110011","111111111111111000","111111111111010110","000000000000010011","111111111111111000","000000000000011001","000000000000001110","111111111111111111","111111111111111111","111111111111101101","111111111111010000","111111111111110100","000000000000011010","111111111111111010","000000000000010011","000000000000001010","000000000000011010","000000000000010110","000000000000000000","000000000000001011","111111111111110111","000000000000001000","111111111111110111","000000000000100110","111111111111111000","000000000000000000","000000000000101100","000000000000011000","000000000000010000","111111111111110011","111111111111111111","111111111111101111","111111111111111100","111111111111111011","000000000000000100","111111111111100101","111111111111100000","000000000000100101","111111111111011111","000000000000000001","000000000000010110","000000000000000010","111111111111111110","000000000000000100","000000000000000010","000000000000000011","111111111111110000","000000000000000100","111111111111101100","000000000000100010","111111111111110101","111111111111111101","000000000000000101","111111111111111110","000000000000000011","000000000000000110","000000000000001001","111111111111111110","000000000000101110","000000000000010011","111111111111111010","000000000000000010","111111111111110010","000000000000001110","000000000000010100","111111111111110001","111111111111111011","111111111111111011","000000000000001111","111111111111111110","000000000000011100","111111111111111110"),
("000000000000010100","111111111111100101","111111111111101100","000000000000000100","000000000000000100","000000000000101001","000000000000010000","000000000000011000","000000000000000101","111111111111100010","000000000000011011","000000000000011011","000000000000010010","111111111111110010","111111111111100100","000000000000001110","000000000000101100","000000000000100001","000000000000010001","000000000000000000","111111111111101011","111111111111011001","111111111111101011","111111111111110000","000000000000000011","000000000000110010","111111111111100110","000000000000000000","111111111111111100","000000000000010000","000000000000100000","111111111111101111","000000000000100110","111111111111111110","000000000000001001","000000000000001010","000000000000000010","000000000000001110","000000000000001110","000000000000000010","111111111111101101","000000000000001010","111111111111110011","111111111111110000","000000000000001111","000000000000000010","111111111111111110","000000000000010000","111111111111111111","111111111111100011","000000000000001101","000000000000101110","111111111111101001","000000000000001000","000000000000001011","111111111111111100","000000000000000111","000000000000000101","111111111111110011","111111111111111101","000000000000010000","111111111111111111","000000000000000011","111111111111101001","111111111111100101","111111111111101001","000000000000001101","000000000000101000","000000000000100111","111111111111100101","000000000000001010","000000000000001010","000000000000000110","000000000000100110","000000000000000011","000000000000101010","000000000000000000","000000000000000110","111111111111100001","000000000000000111","000000000000000100","000000000000001010","000000000000010101","111111111111101010","000000000000101001","111111111111100101","111111111111111110","000000000000001010","000000000000000000","000000000000000000","111111111111110000","000000000000000000","111111111111110010","000000000000001111","111111111111111010","000000000000011100","000000000000000101","000000000000011101","111111111111110000","111111111111000111","000000000000010000","000000000000000110","000000000000010001","000000000000011110","111111111111110110","000000000000101010","000000000000000010","111111111111001010","000000000000000011","111111111111101100","111111111111100111","000000000000010000","000000000000011001","111111111111111100","111111111111011111","000000000000011101","000000000000000010","000000000000010000","111111111111110001","000000000000011100","000000000000001100","000000000000010010","111111111111100100","111111111111000111","111111111111101011","111111111111101110","111111111111111110","000000000000001101"),
("000000000000001010","111111111111001111","111111111111111011","000000000000000111","000000000000010101","000000000000100100","000000000000001000","000000000000010001","000000000000011101","111111111111001111","000000000000001101","000000000000000111","000000000000001010","111111111111101110","111111111111010010","000000000000001100","000000000000000000","000000000000000110","000000000000011010","111111111111111111","000000000000000000","111111111111101001","111111111111111001","111111111111100101","111111111111101100","000000000000011011","111111111111110101","000000000000010011","111111111111111111","000000000000010011","000000000000011000","000000000000000111","111111111111110100","111111111111110111","000000000000000101","000000000000010000","111111111111110100","000000000000000001","000000000000101000","111111111111111100","000000000000011000","111111111111111010","000000000000000010","111111111111011001","111111111111110010","000000000000000111","000000000000010001","111111111111110111","111111111111111010","000000000000000001","000000000000000111","111111111111111100","000000000000001001","000000000000100000","000000000000000100","111111111111101111","111111111111111001","111111111111101000","000000000000000010","000000000000001111","000000000000000101","000000000000000010","111111111111101001","111111111111011100","000000000000000000","000000000000000110","000000000000000010","111111111111110010","000000000000011100","111111111111111001","000000000000001010","000000000000010100","111111111111111010","111111111111111100","000000000000011001","000000000000000000","000000000000010000","111111111111110101","111111111111011010","000000000000000100","000000000000001010","111111111111111111","111111111111111001","000000000000000010","000000000000001010","111111111111101110","111111111111100011","111111111111111011","111111111111111100","000000000000011000","111111111111111000","111111111111110011","111111111111101010","111111111111101000","111111111111101110","000000000000010101","000000000000001000","000000000000001000","111111111111011011","000000000000010010","000000000000010100","000000000000000001","111111111111100100","000000000000010111","111111111111100100","111111111111110110","111111111111111111","000000000000000011","000000000000110101","111111111111110101","000000000000010011","000000000000000100","000000000000001111","000000000000000100","000000000000000110","111111111111110001","111111111111111100","111111111111110110","000000000000011100","000000000000000000","000000000000000101","111111111111111101","000000000000001101","111111111111011110","111111111111110011","000000000000000010","111111111111111100","000000000000010100"),
("111111111111111110","111111111111000001","111111111110111110","000000000000001001","000000000000011100","000000000000011010","000000000000000010","000000000000010001","000000000000000010","111111111111001001","000000000000010011","111111111111111000","000000000000101101","000000000000000000","111111111111010100","000000000000001000","111111111111111001","000000000000101100","000000000000100100","111111111111110110","000000000000000111","000000000000111010","000000000000011010","111111111111110101","111111111111101010","111111111111111001","000000000000000001","111111111111111110","000000000000000011","000000000000011101","000000000000010000","111111111111110100","111111111111101011","111111111111101111","111111111111111010","000000000000001100","111111111111110011","000000000000000101","000000000000110000","111111111111100011","000000000000000111","000000000000000010","111111111111111110","111111111111101100","111111111111011001","000000000000000000","000000000000001001","000000000000010010","111111111111100110","000000000000001001","000000000000011110","111111111111101110","000000000000000110","000000000000100011","000000000000001101","111111111111111000","000000000000001010","111111111111101100","000000000000001101","111111111111111100","000000000000000110","000000000000010111","000000000000001000","111111111111110110","111111111111010110","000000000000000010","111111111111111010","000000000000001010","000000000000010100","111111111111101010","000000000000010110","000000000000001001","111111111111011000","111111111111101110","000000000000010011","000000000000001010","111111111111110101","111111111111101000","111111111111100011","000000000000000110","111111111111111100","111111111111100100","000000000000011001","000000000000010011","000000000000001010","111111111111101001","111111111111100100","111111111111100100","111111111111111100","000000000000000101","000000000000000011","111111111111100101","111111111111011011","000000000000001010","111111111111110101","000000000000011011","111111111111100110","111111111111110100","111111111111011110","000000000000000011","000000000000000000","111111111111110010","111111111111111101","000000000000011111","111111111111111110","000000000000100010","111111111111111000","000000000000001000","000000000000100001","111111111111110000","111111111111110100","000000000000011011","111111111111011100","000000000000001110","000000000000001100","000000000000001001","111111111111110110","000000000000011010","000000000000001111","000000000000000110","000000000000011000","111111111111111110","111111111111100101","111111111111101010","111111111111111110","111111111111110101","111111111111111110","000000000000001010"),
("111111111111111101","111111111111100000","111111111111001000","000000000000100100","000000000000001111","111111111111101111","000000000000001101","000000000000011000","000000000000100110","111111111111100001","000000000000100011","111111111111111111","000000000000011101","000000000000000111","111111111111001111","000000000000011010","111111111111101110","000000000000011100","000000000000000101","000000000000000101","000000000000011101","000000000000110101","000000000000011010","000000000000000001","000000000000001010","111111111111110100","000000000000010000","111111111111111111","111111111111110110","111111111111111110","000000000000000000","000000000000000000","000000000000000011","111111111111101010","111111111111101111","000000000000010000","111111111111100101","000000000000010101","000000000000011101","111111111111100110","000000000000011110","111111111111100100","111111111111101110","111111111111011110","000000000000000000","111111111111110011","000000000000000001","111111111111101001","111111111111110101","111111111111110111","000000000000001110","000000000000000010","000000000000011111","000000000000010000","111111111111111011","111111111111110100","111111111111101011","000000000000010100","000000000000000110","111111111111110101","111111111111110111","111111111111111001","111111111111111100","000000000000010001","111111111111000001","111111111111100111","000000000000011010","111111111111111110","000000000000001001","000000000000010000","000000000000001011","000000000000011010","111111111111100111","111111111111101110","000000000000010001","000000000000001001","111111111111111011","111111111111111111","111111111111111011","000000000000010110","111111111111100111","111111111111111100","111111111111111001","000000000000000001","000000000000010111","111111111111110010","000000000000000000","111111111111111010","111111111111110001","111111111111110110","000000000000000001","111111111111111111","111111111111100111","000000000000000001","111111111111010101","000000000000011110","000000000000000100","111111111111100111","111111111110110100","111111111111100111","000000000000000010","111111111111101110","000000000000000100","000000000000001101","111111111111111001","000000000000101111","111111111111111001","111111111111111101","000000000000111110","111111111111100111","000000000000001000","000000000000000000","111111111111110011","000000000000010011","111111111111111101","000000000000001000","111111111111100110","000000000000000000","000000000000010111","000000000000011110","000000000000001110","000000000000010101","111111111111001101","000000000000000011","111111111111100111","111111111111111000","000000000000001001","111111111111110100"),
("111111111111011010","111111111111011101","111111111111001101","000000000000011011","111111111111111110","111111111111110000","000000000000001011","000000000000010001","000000000000100011","000000000000000111","000000000000000111","111111111111110100","000000000000100000","000000000000000001","111111111111001110","000000000000000011","111111111111110110","000000000000101010","000000000000001111","000000000000000100","111111111111101100","000000000001000000","000000000000010100","111111111111111100","000000000000001000","000000000000010111","000000000000001010","111111111111110110","000000000000010101","000000000000000100","000000000000000000","000000000000000010","000000000000010000","111111111111101010","000000000000001010","000000000000010011","000000000000000110","000000000000001111","000000000000100000","111111111111101000","000000000000001001","000000000000001010","111111111111011101","111111111111011010","111111111111100111","111111111111101000","111111111111100010","000000000000001101","111111111111111100","111111111111101111","000000000000010101","000000000000000000","000000000000100001","000000000000010000","000000000000010000","111111111111110011","111111111111110011","111111111111110101","000000000000011010","111111111111111000","111111111111110001","111111111111110000","111111111111110010","111111111111110101","111111111110111011","000000000000001011","000000000000001001","111111111111111110","111111111111101111","111111111111111010","000000000000010001","111111111111111111","111111111111100100","000000000000000010","000000000000010010","000000000000001000","111111111111110011","000000000000001111","000000000000001001","111111111111111011","111111111111101100","111111111111101000","111111111111110100","000000000000010100","000000000000101001","111111111111111100","111111111111111101","000000000000000000","111111111111101111","111111111111111101","111111111111111100","111111111111111001","111111111111100110","111111111111110110","111111111111101011","000000000000100001","111111111111111010","111111111111110001","111111111111010100","000000000000000000","000000000000000010","111111111111111101","000000000000011000","000000000000010011","000000000000001111","000000000000100110","000000000000010010","000000000000000101","000000000000010100","111111111111111101","000000000000001011","000000000000000111","111111111111101011","111111111111110100","000000000000001001","111111111111111110","111111111111111011","000000000000001111","000000000000000011","000000000000000011","000000000000001011","000000000000000111","111111111111010100","111111111111111001","111111111111111100","111111111111101111","000000000000001100","000000000000000010"),
("111111111111100110","111111111111001010","111111111111011000","000000000000100000","000000000000011011","000000000000001100","000000000000101101","111111111111110000","000000000000000100","000000000000000000","000000000000011111","111111111111110011","000000000000010010","111111111111110010","111111111111010001","000000000000010011","111111111111101100","000000000000001111","000000000000000100","111111111111110111","000000000000000011","000000000001001010","000000000000100000","111111111111111101","111111111111111010","111111111111111011","000000000000000000","111111111111101111","000000000000000011","000000000000011000","000000000000000000","111111111111101110","000000000000000010","111111111111110101","000000000000001000","111111111111101111","000000000000010000","111111111111110011","000000000000011010","111111111111110001","000000000000101100","111111111111111000","111111111111100001","111111111111101101","111111111111111010","111111111111100111","111111111111011010","111111111111111101","111111111111100011","000000000000000111","000000000000010011","111111111111111111","000000000000000011","000000000000100100","000000000000000010","111111111111111110","111111111111100111","000000000000000111","000000000000001100","111111111111111100","000000000000001000","000000000000000111","111111111111110101","000000000000000010","000000000000000110","000000000000001010","000000000000000101","000000000000010100","000000000000000000","111111111111111010","000000000000001001","000000000000010000","000000000000000101","111111111111100001","111111111111110111","000000000000100111","000000000000010001","000000000000001111","000000000000010100","000000000000001000","000000000000000011","111111111111011101","111111111111111010","111111111111101000","000000000000100110","111111111111101101","000000000000001011","000000000000001100","111111111111110101","111111111111111101","000000000000000111","000000000000000101","111111111111111110","000000000000001001","111111111111101010","000000000000100011","000000000000001100","111111111111101100","111111111111100011","111111111111111000","111111111111101111","111111111111100000","000000000000010011","000000000000010011","111111111111110010","000000000000100001","111111111111110000","111111111111101100","000000000000100110","000000000000000011","111111111111101110","000000000000011101","111111111111100111","111111111111110001","000000000000000000","000000000000100111","111111111111111010","000000000000000100","000000000000000000","000000000000010000","111111111111110011","000000000000000101","000000000000010110","111111111111101110","111111111111100100","111111111111100111","111111111111111111","111111111111111000"),
("111111111111101001","111111111111001001","111111111111101011","000000000000001111","000000000000011001","111111111111101100","000000000000110001","111111111111110100","000000000000010000","111111111111111101","000000000000100101","111111111111111010","000000000000000011","111111111111101000","111111111111100111","000000000000100100","111111111111100101","000000000000000100","111111111111101001","000000000000001110","111111111111110010","000000000000010010","000000000000001000","111111111111111000","000000000000000000","000000000000001001","000000000000001001","000000000000000000","111111111111101101","000000000000000100","000000000000001000","000000000000000110","111111111111111100","111111111111101110","000000000000001011","000000000000001111","000000000000000111","111111111111111100","000000000000001000","111111111111011001","000000000000010100","111111111111111100","111111111111011111","000000000000000110","111111111111100010","111111111111101010","111111111111111110","000000000000001110","111111111111101000","000000000000000100","000000000000010001","000000000000001110","000000000000001000","000000000000001001","000000000000010101","111111111111110100","111111111111101101","111111111111110110","000000000000010111","000000000000000000","000000000000001001","111111111111101010","111111111111111100","000000000000000111","000000000000000000","000000000000010111","000000000000100011","000000000000010101","111111111111011100","000000000000010011","111111111111111101","000000000000001010","000000000000010101","111111111111111011","111111111111111111","000000000000100101","111111111111111011","000000000000001011","000000000000010001","000000000000000000","111111111111110101","111111111111100011","111111111111100100","111111111111101010","000000000000010111","111111111111110010","000000000000001110","000000000000000011","111111111111100110","000000000000000011","111111111111111110","111111111111111010","000000000000010010","111111111111111000","111111111111101110","000000000000011011","000000000000001010","111111111111110001","111111111111100101","111111111111111001","000000000000000110","000000000000000011","000000000000000011","000000000000001001","000000000000010011","000000000000000101","111111111111111011","000000000000000101","000000000000100100","000000000000001010","111111111111111100","000000000000101111","111111111111110000","111111111111110111","111111111111100100","000000000000010101","111111111111110111","000000000000100100","000000000000010000","000000000000011100","000000000000010100","000000000000000101","000000000000100001","000000000000000010","111111111111101111","111111111111111110","000000000000001100","111111111111011101"),
("111111111111101110","111111111111011010","111111111111101011","000000000000001000","000000000000010001","000000000000001110","000000000000101110","111111111111101001","000000000000010110","111111111111101110","000000000000010110","111111111111100000","000000000000001100","000000000000001101","111111111111110001","000000000000001011","111111111111110111","000000000000011001","111111111111101011","000000000000001110","111111111111010110","111111111111110001","111111111111111010","000000000000001011","000000000000000100","000000000000011001","000000000000010000","000000000000001001","000000000000000010","000000000000100101","111111111111101010","111111111111111111","111111111111111110","000000000000011001","000000000000001001","000000000000001101","111111111111111110","111111111111111101","111111111111111101","111111111111111100","000000000000001101","111111111111111111","111111111111010101","000000000000010110","000000000000000111","000000000000000110","111111111111110100","000000000000001110","000000000000000101","111111111111110010","000000000000000011","000000000000010001","000000000000010111","000000000000001110","000000000000000111","111111111111110110","111111111111101110","111111111111110100","000000000000001111","111111111111101100","000000000000001001","000000000000000000","000000000000010110","000000000000001101","000000000000011101","000000000000011001","000000000000001111","000000000000101101","111111111111111000","000000000000100110","000000000000000101","111111111111111010","111111111111111000","111111111111110010","111111111111111000","000000000000011101","000000000000000000","000000000000011100","000000000000010111","000000000000001010","111111111111111110","111111111111111100","111111111111011001","111111111111110000","111111111111111111","000000000000000000","111111111111111100","111111111111111011","111111111111111111","111111111111101111","111111111111100100","000000000000011010","111111111111110100","111111111111111111","111111111111110000","000000000000010101","000000000000100100","000000000000001101","000000000000000101","000000000000011000","000000000000011011","000000000000001010","000000000000000110","111111111111111001","000000000000010001","000000000000011010","111111111111101000","111111111111110110","000000000000001111","000000000000010101","000000000000000010","000000000000011100","000000000000100011","000000000000000010","111111111111110111","000000000000011100","111111111111111100","000000000000001101","000000000000011110","000000000000001000","000000000000000110","000000000000011110","111111111111110010","111111111111110011","111111111111100111","000000000000100010","000000000000001110","000000000000000000"),
("000000000000000001","111111111111111011","111111111111111111","000000000000010011","000000000000000000","111111111111111101","000000000000001000","111111111111100111","000000000000010001","000000000000000001","000000000000011010","111111111111110101","111111111111011101","111111111111100001","111111111111101001","000000000000110001","111111111111111010","000000000000001001","000000000000010111","000000000000000000","111111111111110110","111111111111001001","000000000000011001","000000000000100000","000000000000000000","000000000000001110","111111111111111011","111111111111110011","111111111111110110","000000000000001100","000000000000000000","111111111111111110","000000000000000111","111111111111110111","000000000000001001","000000000000010001","000000000000010001","111111111111101001","000000000000000010","111111111111111011","000000000000010000","111111111111111010","111111111111101110","111111111111110000","000000000000101001","111111111111111111","000000000000000110","111111111111110001","000000000000010101","111111111111111110","111111111111111100","000000000000100010","000000000000000111","000000000000001010","000000000000010000","111111111111101110","000000000000000010","000000000000001010","111111111111111001","111111111111110111","000000000000010001","111111111111111000","000000000000001110","000000000000010001","111111111111101100","000000000000011011","000000000000100100","000000000000010110","000000000000000111","000000000000100010","000000000000000101","111111111111101110","111111111111100011","000000000000000010","000000000000001011","000000000000101000","000000000000001011","000000000000011000","000000000000000000","000000000000100001","000000000000000011","000000000000000001","111111111111111000","111111111111111010","000000000000010110","111111111111110101","000000000000001110","111111111111111000","111111111111101010","111111111111100001","000000000000000110","000000000000000010","111111111111111000","000000000000000011","111111111111101100","000000000000010111","000000000000010001","111111111111101110","000000000000000000","000000000000010100","111111111111111001","111111111111111011","000000000000101101","000000000000001100","000000000000010001","000000000000010010","111111111111101011","111111111111110100","000000000000001110","111111111111111100","111111111111101011","000000000000110110","000000000000001101","000000000000001110","111111111111101101","000000000000000011","000000000000100001","000000000000000111","000000000000000110","000000000000000000","000000000000000010","000000000000001100","111111111111111011","111111111111101100","111111111111100101","000000000000001100","000000000000010010","111111111111110101"),
("111111111111111001","000000000000000110","000000000000010111","000000000000001101","111111111111110110","000000000000010000","000000000000001000","111111111111111110","111111111111111101","000000000000001111","111111111111110001","111111111111101101","111111111111101010","111111111111101110","000000000000001101","000000000000101010","111111111111110000","000000000000010000","000000000000001011","111111111111110010","000000000000000101","111111111111100010","111111111111110110","000000000000000110","111111111111110111","111111111111111110","000000000000001010","000000000000000100","111111111111011000","000000000000110100","111111111111101100","111111111111101001","000000000000000000","111111111111111110","111111111111111010","000000000000001010","000000000000010101","111111111111111110","111111111111011101","111111111111110110","000000000000000011","000000000000000010","111111111111101100","000000000000001100","000000000000010100","111111111111110011","000000000000001111","111111111111101110","111111111111110110","000000000000010101","111111111111111001","111111111111110011","111111111111110111","000000000000000000","000000000000001011","000000000000000001","111111111111100111","000000000000001010","000000000000011101","111111111111111101","000000000000000100","111111111111100110","111111111111111011","111111111111111001","111111111111100011","000000000000001110","000000000000101011","000000000000011101","000000000000001000","000000000000011000","000000000000001001","111111111111111101","000000000000001010","111111111111101011","111111111111101001","000000000000001111","000000000000011101","000000000000010001","111111111111111001","111111111111110111","111111111111101101","000000000000011000","111111111111011110","000000000000000110","111111111111101101","111111111111101111","111111111111111110","000000000000000000","000000000000010100","111111111111111011","111111111111101110","000000000000010110","000000000000000101","000000000000000101","000000000000001000","000000000000011000","111111111111110111","111111111111111100","111111111111111011","000000000000011100","111111111111111101","000000000000010010","000000000000011101","000000000000011000","000000000000010111","000000000000010000","111111111111111010","000000000000000110","111111111111101001","000000000000010001","111111111111111000","000000000000100100","000000000000001111","111111111111111000","111111111111110000","000000000000001101","000000000000000101","000000000000101001","000000000000001111","000000000000011100","000000000000010101","111111111111110000","111111111111110000","000000000000001000","111111111111110011","000000000000011101","000000000000100110","111111111111111101"),
("000000000000010100","000000000000001000","111111111111111000","000000000000010110","000000000000010001","000000000000010100","111111111111110001","111111111111110100","000000000000000000","000000000000000100","111111111111110110","000000000000000100","111111111111100110","111111111111011000","111111111111111110","000000000000001111","000000000000000110","000000000000011100","111111111111111111","000000000000001101","111111111111111111","111111111111011101","111111111111111011","000000000000010110","111111111111110101","000000000000000111","111111111111111011","000000000000010001","111111111111111011","000000000000000100","111111111111111110","111111111111111000","000000000000000000","000000000000010100","000000000000001111","000000000000010100","111111111111101111","111111111111100101","111111111111101001","111111111111111111","000000000000010001","000000000000000011","000000000000010111","000000000000000011","000000000000010011","000000000000000001","111111111111111110","000000000000001001","000000000000000101","111111111111110110","000000000000000000","000000000000000000","111111111111101111","111111111111101110","111111111111110001","111111111111011111","111111111111101010","111111111111111011","111111111111110010","000000000000000110","000000000000100001","111111111111110001","000000000000000000","000000000000000011","111111111111101110","000000000000011100","000000000000101101","000000000000100011","111111111111100000","111111111111110110","000000000000000101","111111111111110101","111111111111101101","000000000000001111","000000000000001001","000000000000000000","111111111111110100","000000000000001110","111111111111101111","000000000000000000","111111111111111111","000000000000011000","111111111111100111","000000000000010000","000000000000011000","111111111111111000","000000000000011100","000000000000000101","000000000000000001","000000000000000100","111111111111111001","000000000000011000","111111111111110111","000000000000011001","000000000000000110","000000000000000000","000000000000000000","000000000000000000","111111111111111111","000000000000000100","111111111111110000","000000000000000000","000000000000010110","000000000000010101","000000000000011101","111111111111111110","111111111111111010","000000000000000110","111111111111100101","000000000000000000","111111111111110010","000000000000011100","000000000000011110","111111111111110101","111111111111110011","000000000000011000","000000000000010110","000000000000011000","111111111111101011","000000000000001101","000000000000001111","111111111111100101","000000000000001010","000000000000010111","111111111111001001","000000000000100010","000000000000010100","111111111111111011"),
("000000000000100001","000000000000000100","000000000000010011","000000000000000010","111111111111111011","111111111111111010","111111111111011101","111111111111101011","111111111111111111","000000000000000011","000000000000011011","000000000000001110","111111111111110011","111111111111100101","111111111111111110","000000000000010111","111111111111111111","000000000000010000","000000000000010010","000000000000000110","000000000000011001","111111111111011001","000000000000001110","000000000000001100","111111111111110101","111111111111111010","111111111111111001","000000000000001100","000000000000000001","000000000000100010","111111111111011111","000000000000000001","000000000000011010","000000000000100100","000000000000001001","111111111111111100","000000000000010101","000000000000010000","111111111111100000","000000000000001010","000000000000000100","111111111111111101","000000000000001100","000000000000001011","111111111111111111","111111111111111110","000000000000000101","111111111111110011","111111111111111010","111111111111111000","111111111111011011","000000000000010100","111111111111101011","000000000000001111","000000000000000000","111111111111101011","000000000000000110","000000000000010111","000000000000001000","111111111111110000","000000000000001110","000000000000000110","111111111111100111","000000000000001011","000000000000000001","000000000000011000","000000000000010001","000000000000011001","000000000000000011","111111111111110100","000000000000000111","000000000000000111","111111111111100000","000000000000000110","000000000000000100","000000000000000110","111111111111110011","000000000000000011","000000000000000111","111111111111101110","000000000000010101","000000000000010100","111111111111011110","000000000000010000","000000000000000111","111111111111011011","000000000000100000","111111111111101100","000000000000010100","111111111111101011","000000000000010111","000000000000001000","000000000000000010","000000000000010011","000000000000010110","111111111111111010","000000000000010100","111111111111101111","111111111111101111","111111111111111011","111111111111101000","000000000000010001","000000000000100110","000000000000001110","000000000000000001","000000000000010011","000000000000001100","111111111111110001","111111111111100010","000000000000001110","000000000000010011","000000000000100010","000000000000000100","000000000000000000","111111111111111101","000000000000000011","000000000000010001","000000000000011001","000000000000000101","000000000000001001","000000000000001110","111111111111111001","000000000000001110","000000000000001011","111111111111001010","000000000000001100","000000000000000010","000000000000000001"),
("000000000000000101","000000000000000101","111111111111111000","111111111111111100","111111111111111010","111111111111110010","111111111111011000","111111111111101101","111111111111101100","000000000000000111","000000000000001001","000000000000001111","111111111111110101","111111111111011010","111111111111110111","111111111111111011","000000000000010010","111111111111110010","000000000000001110","000000000000011000","000000000000000000","000000000000000011","000000000000100011","111111111111110001","000000000000001111","000000000000000101","000000000000000110","000000000000000100","111111111111111010","000000000000100111","111111111111100110","111111111111111101","111111111111111010","000000000000100001","000000000000000001","000000000000011110","111111111111111110","111111111111101110","000000000000001000","111111111111111100","000000000000001010","000000000000010010","000000000000010011","000000000000010110","000000000000000000","111111111111111010","111111111111110111","111111111111100101","000000000000010100","111111111111111101","111111111111011101","000000000000010001","000000000000000100","111111111111101011","111111111111110111","111111111111110111","000000000000010011","000000000000010011","000000000000001101","111111111111110011","000000000000010000","000000000000000111","111111111111101110","111111111111101010","111111111111110010","000000000000000011","111111111111101111","000000000000001000","111111111111111000","000000000000000111","000000000000010010","000000000000000111","111111111111110010","000000000000001101","000000000000010010","111111111111100101","000000000000001010","000000000000000010","111111111111111010","000000000000001100","000000000000000000","000000000000001100","111111111111010101","111111111111111101","000000000000001001","111111111111110010","000000000000010011","111111111111110100","000000000000010101","000000000000001110","000000000000001001","000000000000100100","000000000000010100","000000000000000100","111111111111110011","111111111111100111","000000000000001011","000000000000000110","000000000000010011","111111111111100010","000000000000000010","000000000000000001","000000000000010011","111111111111111010","000000000000001110","111111111111111010","111111111111111100","111111111111111111","000000000000001000","111111111111101110","111111111111111011","000000000000001100","000000000000001101","111111111111111101","000000000000001011","000000000000000010","000000000000000000","000000000000001100","111111111111110101","000000000000001111","000000000000011011","111111111111100001","000000000000000000","000000000000110000","111111111111011010","000000000000101000","000000000000001000","111111111111110111"),
("000000000000011101","000000000000010101","111111111111101110","000000000000000100","111111111111111110","000000000000000011","111111111111100111","000000000000001001","000000000000000010","111111111111111000","000000000000010011","000000000000101001","111111111111111000","111111111111011100","000000000000011000","000000000000010110","111111111111110011","000000000000001010","111111111111101110","111111111111110001","111111111111111011","000000000000011100","000000000000001001","111111111111100010","000000000000001010","000000000000001111","000000000000001111","000000000000001001","000000000000010010","000000000000100101","000000000000000110","111111111111110101","000000000000010001","000000000000010100","111111111111111010","000000000000000000","000000000000001110","000000000000000000","000000000000001101","000000000000000110","000000000000010010","000000000000010100","111111111111110110","000000000000000010","000000000000010000","111111111111111001","000000000000000101","111111111111011101","000000000000000101","000000000000001110","111111111111110001","000000000000001011","111111111111101010","000000000000001100","111111111111110101","111111111111101000","000000000000010010","000000000000001110","000000000000000011","000000000000010000","000000000000001011","000000000000011001","111111111111100011","111111111111111010","111111111111111100","000000000000001011","111111111111011111","000000000000001110","000000000000010100","111111111111110000","000000000000010010","000000000000001001","111111111111010110","111111111111111011","000000000000001000","111111111111101000","000000000000000100","000000000000001000","111111111111111100","000000000000000100","111111111111111111","000000000000011000","111111111111001011","000000000000010011","000000000000001111","000000000000000101","000000000000010010","111111111111110010","000000000000101101","000000000000010011","000000000000001101","000000000000000000","000000000000100101","111111111111111001","000000000000001110","111111111111011111","000000000000001110","111111111111101110","000000000000001001","111111111111101100","111111111111110010","000000000000001101","000000000000010010","000000000000001001","111111111111101000","000000000000000000","000000000000000010","111111111111101111","000000000000010011","111111111111111110","111111111111110101","000000000000101111","000000000000001110","000000000000001110","111111111111111000","111111111111111110","000000000000000001","111111111111110011","111111111111110011","000000000000010110","000000000000001101","000000000000000111","111111111111101000","000000000000100010","111111111111010111","000000000000010001","000000000000000110","111111111111110011"),
("000000000000011010","000000000000101010","000000000000000101","000000000000001110","111111111111111110","000000000000001001","111111111111101110","111111111111101101","111111111111110101","000000000000000110","000000000000100111","000000000000100110","111111111111110011","111111111111101010","111111111111101110","000000000000011101","000000000000000110","000000000000010010","111111111111111110","000000000000000100","000000000000010010","000000000000100001","000000000000011101","111111111111110100","000000000000001000","111111111111111001","000000000000001000","111111111111111111","111111111111110101","000000000000001000","000000000000010001","111111111111111111","111111111111110010","111111111111111111","111111111111101001","000000000000010001","000000000000000011","000000000000010011","000000000000011001","000000000000000000","000000000000001011","000000000000010010","111111111111110001","000000000000000000","000000000000011111","111111111111110111","111111111111100011","111111111111101101","000000000000001001","000000000000001010","111111111111101000","000000000000010010","111111111111111111","000000000000000001","000000000000001011","000000000000000010","000000000000010001","000000000000000100","111111111111100100","111111111111111000","111111111111101101","000000000000010010","111111111111101100","111111111111110001","111111111111110011","000000000000000011","111111111110111010","111111111111111101","111111111111110110","111111111111110000","000000000000011000","000000000000001000","111111111111111010","111111111111110010","000000000000011000","111111111111010010","111111111111110101","111111111111111011","111111111111110000","111111111111111001","000000000000001011","000000000000000011","111111111111010111","111111111111100111","000000000000011000","111111111111101010","111111111111111000","000000000000001010","000000000000010011","000000000000001111","111111111111111110","000000000000010000","000000000000100000","111111111111111100","111111111111110011","111111111111011100","000000000000001101","000000000000000001","111111111111110001","111111111111100100","111111111111110101","111111111111111100","000000000000000000","000000000000011100","111111111111101110","111111111111111110","111111111111111011","111111111111011001","111111111111110001","111111111111101110","111111111111111110","000000000000000100","000000000000010100","000000000000000100","111111111111110100","000000000000000100","000000000000011000","000000000000011000","000000000000001101","000000000000010011","000000000000010001","111111111111100101","000000000000001100","000000000000001110","111111111111010010","000000000000001001","000000000000011000","000000000000000110"),
("000000000000000101","000000000000011000","111111111111110000","000000000000011011","000000000000000011","000000000000010101","111111111111101011","000000000000000100","000000000000001100","000000000000000011","000000000000110000","000000000000011110","000000000000000101","111111111111100000","111111111111100110","000000000000100011","000000000000000100","000000000000010000","000000000000001111","000000000000001110","111111111111110000","000000000000011010","000000000000000000","111111111111101110","000000000000000010","000000000000010011","000000000000011011","000000000000001101","111111111111111110","000000000000001011","000000000000011111","111111111111100110","000000000000000000","111111111111111010","000000000000010000","111111111111111111","111111111111011101","111111111111110110","000000000000011000","000000000000010100","000000000000011100","111111111111110110","000000000000001001","000000000000000001","000000000000011000","111111111111110110","000000000000000010","111111111111110010","000000000000000001","111111111111011110","111111111111100011","111111111111111011","111111111111110111","111111111111111001","111111111111111101","000000000000000000","111111111111110110","000000000000001100","111111111111110110","111111111111111000","111111111111100001","000000000000010111","111111111111101001","000000000000001010","000000000000010001","000000000000000011","111111111110110000","111111111111111110","000000000000000011","000000000000010000","000000000000000001","000000000000100100","111111111111111111","111111111111111101","000000000000001110","111111111111100100","111111111111110100","000000000000001010","000000000000000000","111111111111100010","000000000000011001","000000000000000000","111111111111010010","111111111111001100","000000000000001101","111111111111101001","111111111111111100","000000000000000000","000000000000011000","000000000000011110","000000000000001101","000000000000000100","000000000000000101","111111111111101101","000000000000000001","111111111111010000","111111111111110101","111111111111110101","111111111111110001","111111111111111010","000000000000001111","000000000000000000","111111111111110101","000000000000011101","111111111111101001","111111111111111011","000000000000001010","111111111111110011","000000000000000101","111111111111100010","000000000000001101","000000000000011101","000000000000000000","000000000000000111","111111111111110000","111111111111111000","111111111111110110","000000000000001001","111111111111100000","111111111111111010","000000000000010101","111111111111101100","000000000000000110","000000000000001010","111111111111011001","000000000000001001","000000000000011100","000000000000001100"),
("000000000000000000","000000000000101111","111111111111100010","000000000000000000","000000000000001010","000000000000011111","111111111111110000","000000000000011100","111111111111110010","000000000000000110","000000000000010110","000000000000110101","111111111111101001","111111111111010111","000000000000000010","000000000000010111","000000000000011001","000000000000000011","000000000000000000","000000000000010011","111111111111100100","000000000000000000","000000000000000101","111111111111010100","111111111111101100","000000000000010011","000000000000000100","000000000000001000","000000000000001101","111111111111111000","111111111111110110","111111111111100011","111111111111110100","000000000000000101","000000000000011011","000000000000011111","111111111111100101","000000000000011011","000000000000000000","000000000000100001","000000000000000010","111111111111101011","111111111111110010","111111111111111011","000000000000000000","111111111111110111","111111111111110100","000000000000010100","000000000000000001","111111111111101011","111111111111101010","000000000000000000","111111111111100001","000000000000000111","111111111111111110","111111111111101110","111111111111011110","111111111111111111","111111111111110100","000000000000000000","111111111111100011","000000000000001011","000000000000010000","000000000000001000","111111111111110000","111111111111110101","111111111110101000","000000000000001110","111111111111101111","111111111111111111","000000000000000000","000000000000010010","111111111111001100","000000000000000001","000000000000101101","111111111111010111","000000000000001001","000000000000010000","111111111111011101","000000000000001000","111111111111101111","111111111111111000","111111111111100010","111111111111010111","000000000000001101","111111111111111111","111111111111110010","111111111111111111","111111111111111110","000000000000010100","000000000000011001","111111111111100101","111111111111101010","111111111111011100","111111111111011011","111111111111010000","111111111111101010","111111111111101010","111111111111010000","111111111111111101","000000000000000001","000000000000001110","111111111111001110","000000000000010111","000000000000000111","111111111111100100","111111111111111010","111111111111010110","111111111111110111","111111111111100001","000000000000000010","000000000000001000","000000000000010000","111111111111111000","111111111111110010","111111111111110111","111111111111101100","000000000000001101","111111111111101010","000000000000011011","000000000000011001","000000000000010000","111111111111110110","000000000000001010","111111111111111000","000000000000001100","000000000000010111","111111111111111010"),
("000000000000001110","000000000000011000","000000000000001010","111111111111111101","000000000000100010","000000000000100010","111111111111011011","000000000000001000","111111111111110101","000000000000000001","000000000000010100","000000000000101010","000000000000000010","000000000000010010","111111111111110001","111111111111111011","000000000000010001","111111111111101111","111111111111100000","111111111111110100","000000000000000011","111111111111110000","000000000000011000","111111111111100011","111111111111101000","000000000000011010","000000000000011011","000000000000100000","111111111111111000","000000000000000001","000000000000010110","111111111111111100","111111111111010101","111111111111111100","000000000000000111","000000000000000110","111111111111110111","000000000000001001","000000000000001011","111111111111101110","000000000000010010","000000000000001011","000000000000001001","000000000000010110","000000000000011110","111111111111110110","111111111111100001","000000000000010010","111111111111110101","111111111111100011","000000000000000001","000000000000001111","111111111111010010","000000000000101101","000000000000001010","000000000000010000","111111111111011110","111111111111101101","111111111111110111","000000000000001101","111111111111010110","000000000000010010","000000000000000111","111111111111111101","111111111111101010","111111111111011111","111111111111001010","111111111111100010","111111111111110001","111111111111100110","000000000000001001","000000000000000000","111111111110110001","111111111111110010","000000000000011010","111111111111100000","111111111111110110","111111111111111011","111111111111111101","111111111111101010","111111111111111011","111111111111111100","111111111111110101","111111111111101001","000000000000100011","000000000000000011","111111111111011100","000000000000011001","000000000000000101","000000000000000000","000000000000010010","111111111111110111","000000000000000001","111111111111111010","000000000000000000","111111111111101110","000000000000001011","111111111111011110","111111111111011010","000000000000000111","111111111111111101","111111111111111010","111111111111001011","111111111111111111","111111111111101000","111111111111110000","000000000000000011","111111111111011010","000000000000001111","111111111111011000","111111111111111111","000000000000001101","000000000000001001","000000000000001111","111111111111011111","111111111111100010","111111111111111011","000000000000000011","111111111111010000","000000000000001111","111111111111111001","111111111111111111","000000000000001001","000000000000000010","111111111111010100","000000000000000111","111111111111111010","000000000000001100"),
("000000000000100110","000000000000001000","000000000000000010","000000000000000101","000000000000111011","000000000000110100","000000000000001010","000000000000001101","000000000000001011","000000000000001010","000000000000010100","000000000000000011","000000000000000001","000000000000001011","111111111111001110","000000000000000111","000000000000010000","111111111111111110","111111111111110001","111111111111111000","111111111111110100","111111111111101000","000000000000010111","111111111111101001","111111111111010101","000000000000000110","000000000000010001","000000000000001100","000000000000001101","000000000000000010","000000000000001111","111111111111010001","000000000000000000","111111111111110110","111111111111111000","000000000000000111","111111111111110101","000000000000001101","111111111111100000","111111111111110011","000000000000010000","111111111111111001","000000000000000100","000000000000010101","000000000000101010","111111111111100000","111111111111100010","000000000000000110","111111111111110110","111111111111100000","111111111111010110","000000000000000100","111111111111011000","000000000000011010","111111111111101101","000000000000100100","111111111111000110","111111111111110000","111111111111100110","111111111111111011","111111111111011011","000000000000000110","000000000000000100","000000000000010000","000000000000001010","111111111111111100","111111111111100000","111111111111111001","111111111111110000","111111111111101100","000000000000010010","111111111111101010","111111111111001101","000000000000000110","111111111111111110","111111111111111100","111111111111111111","111111111111101101","111111111111100100","111111111111111111","111111111111111010","000000000000001110","000000000000010000","000000000000000010","000000000000000011","000000000000001101","111111111111011011","111111111111111101","111111111111101100","111111111111011101","111111111111111100","111111111111010110","000000000000000010","111111111111100101","111111111111111101","111111111111010101","111111111111100110","111111111111111101","111111111110111010","000000000000010001","000000000000001011","111111111111111010","111111111110110010","000000000000000110","111111111111101100","111111111111111101","000000000000010100","111111111111010011","111111111111111011","111111111111110100","111111111111111001","000000000000010101","000000000000000011","000000000000001010","000000000000011000","111111111111010010","111111111111011110","000000000000001011","111111111111010011","111111111111101101","111111111111111011","111111111111110010","000000000000000100","000000000000010101","111111111111110010","000000000000000111","111111111111110110","111111111111111100"),
("111111111111101110","000000000000010101","000000000000001111","000000000000011010","000000000000011100","000000000000011011","111111111111111011","000000000000010101","000000000000000000","000000000000000100","000000000000100110","000000000000000111","000000000000000000","000000000000100011","111111111111011110","111111111111111111","000000000000001011","000000000000010000","111111111111101100","000000000000001110","111111111111100101","111111111111001101","000000000000011110","111111111111110110","111111111111111011","000000000000010000","000000000000000101","000000000000010110","111111111111101010","111111111111110001","000000000000001001","111111111111100101","000000000000000111","111111111111111001","111111111111101011","111111111111101110","000000000000000000","000000000000000110","111111111111101101","111111111111111011","111111111111111101","111111111111111011","111111111111101111","111111111111111100","000000000000010010","111111111111110000","111111111111101101","111111111111111111","111111111111101100","000000000000000100","000000000000001010","000000000000100011","111111111111101100","000000000000001011","000000000000001011","000000000000001001","111111111111101110","111111111111110001","111111111111111001","000000000000000101","111111111111000101","000000000000000000","000000000000100101","000000000000011001","111111111111011011","111111111111101001","111111111111111010","111111111111101111","111111111111110110","111111111111110001","000000000000001100","111111111111110010","111111111111100011","000000000000000001","000000000000000000","000000000000000111","111111111111110011","000000000000001111","111111111111101011","000000000000000000","111111111111101011","000000000000101010","000000000000011001","111111111111101010","000000000000000010","111111111111110110","111111111111111001","000000000000001000","000000000000001000","111111111111100100","111111111111011101","111111111111111111","111111111111101110","000000000000001001","111111111111111101","111111111111100000","000000000000011001","000000000000000000","000000000000000011","111111111111110110","000000000000010000","000000000000000000","111111111111001101","000000000000011010","000000000000000001","111111111111110101","111111111111111100","111111111111010100","111111111111100010","111111111111100111","000000000000010010","000000000000011010","111111111111101111","111111111111110111","000000000000010110","111111111111110101","111111111111011010","111111111111111011","111111111111010011","111111111111111110","000000000000001110","111111111111101110","111111111111110101","111111111111110110","111111111111010100","111111111111110000","111111111111110011","000000000000011000"),
("000000000000101000","000000000000011000","000000000000011000","111111111111111110","111111111111110100","111111111111111110","111111111111110001","000000000000001010","111111111111111011","000000000000000111","000000000000010010","111111111111110001","000000000000101101","000000000000011110","111111111111111001","000000000000000000","111111111111111110","000000000000001110","111111111111011110","000000000000000100","000000000000001100","111111111111110000","000000000000000011","000000000000001110","000000000000001000","000000000000001110","000000000000001110","000000000000100011","111111111111011111","000000000000001100","000000000000101001","111111111111010000","000000000000010100","000000000000000000","111111111111111111","111111111111101000","111111111111110001","000000000000001110","000000000000000000","000000000000000010","000000000000011010","111111111111110010","000000000000000010","000000000000000110","000000000000111001","111111111111011101","111111111111011001","111111111111011110","111111111111101101","111111111111101000","111111111111110100","000000000000110000","111111111111101101","000000000000101111","000000000000000011","000000000000101000","111111111111110111","000000000000000011","111111111111100111","000000000000000100","111111111111010010","000000000000011001","111111111111110110","000000000000000000","000000000000010100","111111111111110101","111111111111101001","111111111111101110","111111111111110101","111111111111110010","000000000000010110","000000000000011000","111111111111111001","111111111111110010","111111111111111000","111111111111111011","000000000000101100","111111111111110101","000000000000000100","111111111111110010","111111111111101110","000000000000011011","000000000000000000","111111111111101100","000000000000100111","000000000000000110","000000000000010000","000000000000001101","111111111111110010","111111111111010011","111111111111011010","111111111111101110","000000000000000001","111111111111011011","000000000000001110","000000000000000001","000000000000001010","000000000000100000","000000000000010000","000000000000001011","000000000000000000","111111111111111101","111111111111010101","000000000000000001","111111111111101101","111111111111111000","111111111111111100","111111111111001100","111111111111001100","111111111111110010","000000000000000000","000000000000010001","000000000000000001","111111111111101011","000000000000100000","111111111111011100","111111111111010010","000000000000000100","111111111111110110","000000000000010100","000000000000100001","000000000000001110","000000000000010010","000000000000010011","111111111111011011","111111111111110000","000000000000000100","111111111111100101"),
("000000000000011001","000000000000001011","000000000000110011","000000000000100001","000000000000010110","111111111111110101","111111111111111100","000000000000000110","111111111111100000","111111111111010111","000000000000100011","111111111111101011","000000000000111100","000000000000011111","000000000000010100","000000000000001111","111111111111100101","000000000000100001","111111111111111000","111111111111111000","000000000000010011","000000000000000111","000000000000000010","000000000000010101","111111111111111000","000000000000001111","000000000000000000","000000000000100101","000000000000000100","111111111111101101","000000000001000110","111111111111011011","111111111111111101","111111111111110111","000000000000001001","111111111111011010","000000000000010011","000000000000010100","111111111111101010","000000000000000111","000000000000000111","111111111111100010","111111111111111001","000000000000001011","000000000000000101","111111111111111010","111111111110111111","111111111111111010","111111111111100101","111111111111001100","111111111111001100","000000000000001110","111111111111100000","000000000000011001","000000000000110111","000000000000101111","000000000000000010","111111111111110000","111111111111111110","000000000000001100","111111111111101001","000000000000011000","000000000000011011","111111111111100101","000000000000011101","000000000000001100","111111111111111100","111111111111001001","111111111111111101","111111111111101100","111111111111110000","111111111111101110","111111111111011110","111111111111111100","000000000000010010","111111111111110101","000000000000110001","000000000000011110","000000000000001100","111111111111101011","111111111111110011","000000000000001111","000000000000000000","111111111111101101","000000000000001011","000000000000001110","111111111111111101","000000000000001001","111111111111011100","111111111111011111","111111111111101000","111111111111111000","111111111111110110","111111111111100101","000000000000000010","000000000000000100","111111111111111000","111111111111111100","111111111111111011","111111111111111110","000000000000101000","111111111111011110","111111111111110001","111111111111111111","000000000000001011","111111111111110000","111111111111110101","111111111111010111","111111111111001110","000000000000000011","111111111111111101","000000000000101100","111111111110111111","111111111111001110","111111111111110110","111111111111110000","111111111111010001","111111111111010110","000000000000010000","111111111111100101","000000000000011000","000000000000001000","000000000000011010","000000000000001101","111111111111101101","111111111111111001","000000000000001100","111111111111101001"),
("000000000000000010","111111111111111111","000000000000010011","000000000000000010","000000000000000011","111111111111111111","000000000000001001","000000000000000001","000000000000000111","111111111111011001","000000000000000111","111111111111101110","111111111111111101","000000000000011101","000000000000001110","000000000000000001","111111111111111001","000000000000001011","111111111111111010","111111111111110101","000000000000000111","000000000000010000","111111111111110100","000000000000001100","111111111111110100","000000000000001100","000000000000000110","111111111111101010","111111111111111101","000000000000001010","000000000000100101","111111111111111010","111111111111101011","111111111111111010","000000000000011011","000000000000001101","000000000000011000","000000000000001110","111111111111111001","111111111111110010","111111111111110110","111111111111110100","111111111111111001","111111111111110010","111111111111110111","000000000000000100","000000000000000000","111111111111111100","111111111111101101","111111111111011001","111111111111100011","000000000000001000","000000000000010011","000000000000011001","000000000000101100","000000000000000000","111111111111111111","111111111111101111","000000000000001101","111111111111111011","111111111111101100","000000000000010011","111111111111100110","000000000000000100","000000000000011001","111111111111111011","111111111111011110","111111111111101010","000000000000011011","000000000000000100","000000000000001001","111111111111111000","111111111111101000","111111111111111100","111111111111101111","111111111111101111","111111111111111011","000000000000001011","111111111111110111","111111111111101001","000000000000010000","000000000000001110","111111111111100001","000000000000100101","000000000000010010","000000000000010011","111111111111100010","111111111111101001","111111111111111101","000000000000000101","000000000000000110","111111111111100111","111111111111110101","111111111111100011","000000000000001001","111111111111101001","111111111111100111","111111111111100101","111111111111010110","111111111111111011","111111111111111100","111111111111101101","111111111111110000","111111111111110110","000000000000001100","111111111111100100","000000000000000010","111111111111110101","111111111111111101","000000000000010000","000000000000010100","000000000000000100","111111111111001101","111111111111100011","000000000000000000","111111111111100111","111111111111110001","111111111111010000","111111111111101110","111111111111011011","000000000000001110","111111111111111100","111111111111101111","000000000000110001","111111111111100111","000000000000000110","000000000000000000","111111111111110011"),
("111111111111111111","000000000000100111","111111111111111111","111111111111111001","000000000000101001","111111111111111000","111111111111011100","000000000000001111","111111111111101000","000000000000101101","111111111111110011","000000000000011111","111111111111100101","000000000000011110","111111111111110011","111111111111110101","111111111111101101","111111111111110011","111111111111101100","111111111111110111","111111111111110000","111111111111101110","000000000000000111","000000000000000001","000000000000010101","111111111111101110","000000000000010010","111111111111100010","000000000000010111","000000000000010001","000000000000001101","111111111111110000","111111111111101011","000000000000000010","000000000000010010","000000000000011000","000000000000001111","000000000000100010","000000000000001110","000000000000000101","111111111111101100","000000000000011100","111111111111110100","111111111111110010","111111111111111001","000000000000100010","111111111111110010","000000000000011100","000000000000000110","111111111111001011","000000000000000110","000000000000010101","000000000000000100","000000000000011011","111111111111101101","111111111111011011","111111111111110111","111111111111110101","111111111111101101","111111111111110101","000000000000000111","111111111111111101","111111111111101011","000000000000001001","000000000000101110","000000000000001011","000000000000000000","000000000000000011","000000000000011110","000000000000000001","111111111111100100","000000000000010111","000000000000011010","111111111111101001","000000000000000011","111111111111110101","111111111111110001","111111111111111101","111111111111100000","111111111111101110","000000000000001000","000000000000000001","111111111111111100","000000000000101100","000000000000000001","000000000000100010","000000000000011100","000000000000101100","111111111111011100","000000000000101011","000000000000011010","111111111111100111","000000000000100100","111111111111101010","111111111111001111","111111111111100100","000000000000000000","111111111111011100","000000000000011001","111111111111110010","111111111111101011","000000000000011011","111111111111011111","000000000000001001","000000000000000000","111111111111011011","111111111111101101","111111111111111100","000000000000010000","111111111111110001","111111111111100001","000000000000001000","000000000000000101","111111111111110000","111111111111100111","111111111111100110","111111111111101100","000000000000101001","000000000000001001","111111111111111001","000000000000010010","000000000000010000","111111111111100110","111111111111111100","111111111111100010","000000000000010111","111111111111101010","111111111111101000"),
("000000000000000110","111111111111110100","000000000000000101","000000000000000100","111111111111111001","111111111111111010","111111111111110101","000000000000000100","111111111111110010","000000000000010000","000000000000001100","000000000000000011","111111111111101100","000000000000000000","111111111111101101","000000000000001011","111111111111110000","000000000000000110","111111111111110010","000000000000000001","111111111111110011","111111111111101110","111111111111110000","000000000000000110","111111111111101101","000000000000010001","111111111111101100","000000000000001000","000000000000010010","111111111111111111","111111111111110100","000000000000001001","111111111111101110","000000000000001001","111111111111110111","000000000000001110","111111111111110110","000000000000010010","000000000000001110","000000000000001010","000000000000001100","000000000000001011","000000000000001110","111111111111111001","111111111111111001","000000000000010010","111111111111111100","111111111111110010","000000000000000110","000000000000001100","111111111111101110","000000000000001000","111111111111111010","111111111111101100","000000000000000100","000000000000000111","000000000000000001","000000000000001111","000000000000010100","000000000000001101","000000000000000010","000000000000010101","111111111111111010","000000000000000100","000000000000010001","111111111111111111","111111111111110000","111111111111111101","000000000000010011","000000000000000011","111111111111111010","000000000000000111","000000000000000000","000000000000000111","000000000000000100","111111111111111100","111111111111110001","000000000000010001","111111111111101100","000000000000010011","000000000000001011","111111111111111100","000000000000000111","000000000000000010","111111111111110111","111111111111101110","111111111111110000","111111111111110111","111111111111110100","111111111111101101","111111111111110101","000000000000001011","111111111111111001","111111111111110000","000000000000010100","000000000000010001","111111111111101101","111111111111110101","000000000000001010","111111111111111110","000000000000010011","111111111111101011","000000000000000110","111111111111101101","111111111111111011","000000000000010100","000000000000001110","000000000000010010","000000000000000000","000000000000000000","111111111111101111","000000000000010100","111111111111101100","111111111111110000","000000000000010010","111111111111110111","111111111111111010","000000000000001110","000000000000000011","000000000000000100","111111111111110101","111111111111111000","111111111111111000","111111111111110010","000000000000001100","111111111111110010","000000000000001010","111111111111110101"),
("000000000000001001","000000000000001001","000000000000001101","000000000000000011","111111111111101110","000000000000001101","111111111111110110","000000000000001100","000000000000000101","000000000000010011","111111111111101110","111111111111101101","111111111111111011","000000000000010000","111111111111111110","000000000000001111","000000000000001111","000000000000010010","111111111111111000","000000000000010000","000000000000010011","111111111111110001","000000000000001110","111111111111111111","000000000000000101","000000000000000001","111111111111110001","111111111111101110","000000000000001111","000000000000001000","000000000000010100","000000000000000100","111111111111110001","111111111111111101","000000000000000001","000000000000001001","111111111111101110","111111111111110000","000000000000010100","000000000000001011","111111111111111101","111111111111101110","111111111111110100","000000000000010000","111111111111110100","000000000000001011","000000000000000000","000000000000000010","000000000000001101","000000000000001010","111111111111111001","111111111111101101","111111111111110010","000000000000001001","111111111111110111","111111111111111101","000000000000000001","000000000000001001","000000000000000100","111111111111111011","111111111111111111","111111111111101110","111111111111111000","111111111111110100","000000000000001110","000000000000010001","111111111111110010","000000000000000001","000000000000000100","111111111111110011","000000000000000011","111111111111110010","111111111111101100","111111111111111100","111111111111110011","000000000000000110","111111111111111111","000000000000000000","000000000000001010","000000000000001010","111111111111110100","000000000000010011","111111111111111110","000000000000000111","111111111111111011","000000000000000000","111111111111111000","000000000000000110","000000000000001010","111111111111101110","000000000000000111","000000000000001100","000000000000010000","000000000000001111","111111111111110000","111111111111101110","111111111111111110","111111111111110010","000000000000010100","000000000000000110","000000000000001110","111111111111111001","111111111111111111","000000000000001010","111111111111101111","000000000000000100","111111111111111000","111111111111101110","111111111111111010","000000000000000011","111111111111101101","000000000000001010","111111111111111111","000000000000001111","000000000000000101","000000000000000001","000000000000001111","000000000000000001","111111111111110001","000000000000010000","000000000000000110","111111111111110111","111111111111111011","000000000000010000","000000000000000011","000000000000001011","111111111111110010","000000000000000001"),
("000000000000010011","000000000000001011","000000000000000011","111111111111110110","000000000000000111","000000000000000001","000000000000000111","000000000000000110","000000000000010010","111111111111101111","000000000000000111","111111111111110100","000000000000010001","000000000000001011","000000000000000111","000000000000010001","111111111111110101","000000000000001011","000000000000000000","000000000000010100","000000000000010010","111111111111111010","111111111111111100","000000000000000000","000000000000001100","111111111111111011","000000000000001110","111111111111110010","000000000000000000","111111111111110010","000000000000001111","111111111111101111","111111111111101100","000000000000001101","000000000000001100","000000000000010001","111111111111101110","111111111111111010","000000000000000010","111111111111111100","111111111111101101","111111111111110111","000000000000001100","111111111111101110","111111111111110100","000000000000010000","111111111111110101","111111111111111101","000000000000000000","000000000000000000","000000000000000101","000000000000001110","000000000000001011","111111111111111000","111111111111111000","111111111111101100","000000000000010100","111111111111111100","111111111111110011","111111111111111001","000000000000000101","000000000000000101","111111111111110110","111111111111110101","000000000000001010","000000000000001110","111111111111101110","000000000000001110","111111111111111010","111111111111110000","000000000000000100","000000000000000000","111111111111101111","000000000000001010","000000000000001110","000000000000010001","111111111111111011","111111111111110000","000000000000010010","000000000000000110","111111111111101110","111111111111111110","000000000000000110","000000000000010010","000000000000010010","000000000000000101","111111111111111100","000000000000001010","000000000000010000","000000000000001010","000000000000000111","111111111111110101","111111111111111000","111111111111111011","111111111111110000","000000000000001111","111111111111110111","000000000000010001","111111111111110101","000000000000001010","111111111111110111","000000000000010011","111111111111111100","111111111111111000","111111111111111011","000000000000010010","000000000000000110","111111111111110010","111111111111110111","111111111111110000","000000000000001011","000000000000000010","111111111111110111","111111111111111001","111111111111110111","000000000000001010","111111111111110000","000000000000010000","111111111111110111","111111111111101101","000000000000010100","111111111111111001","111111111111101110","000000000000000111","000000000000000111","000000000000001110","000000000000000000","000000000000001110"),
("111111111111110111","111111111111110110","111111111111101000","000000000000010110","111111111111101101","000000000000001000","111111111111100000","000000000000100001","000000000000010101","111111111111111110","000000000000100010","000000000000011000","111111111111110100","111111111111011101","111111111111101010","000000000000000101","000000000000010101","000000000000000101","111111111111110101","000000000000010110","111111111111111011","111111111111110010","000000000000000100","111111111111100100","111111111111111010","000000000000001111","111111111111111101","111111111111111000","000000000000110011","000000000000011100","111111111111101111","000000000000101011","000000000000001001","111111111111111100","111111111111101101","000000000000100000","111111111111110011","000000000000100100","000000000000000000","000000000000010000","111111111111100010","111111111111101010","111111111111110111","111111111111111001","111111111111111110","111111111111110011","111111111111110101","000000000000000010","000000000000001100","000000000000100010","000000000000011011","000000000000000110","111111111111100001","111111111111111111","000000000000100111","111111111111011111","111111111111010011","000000000000010000","111111111111011110","000000000000010010","000000000000100000","000000000000110111","000000000000001111","111111111111111111","111111111111101001","111111111111111000","111111111111011101","000000000000010000","000000000000100011","111111111111100011","000000000000001111","000000000000100000","000000000000011001","111111111111111101","000000000000011110","000000000000001001","111111111111100110","000000000000000101","111111111111100000","000000000000110000","111111111111110111","000000000000010111","111111111111110110","000000000000000011","000000000000001100","111111111111110010","111111111111100011","000000000000001100","000000000000000011","000000000000001000","111111111111110100","000000000000001010","111111111111011111","111111111111100111","111111111111010110","111111111111110110","000000000000101000","111111111111111000","000000000000000111","111111111111110110","000000000000010100","111111111111111111","000000000000000010","000000000000100010","111111111111111000","000000000000010000","111111111111110101","111111111111110010","000000000000010000","111111111111101110","111111111111010111","111111111111110010","000000000000010101","000000000000010100","000000000000111100","000000000000001010","000000000000001010","000000000000001000","111111111111111110","000000000000011010","111111111111111000","111111111111101010","111111111111110100","111111111111100101","111111111111111110","111111111111110111","111111111111111100","111111111111110101"),
("000000000000010001","111111111111101100","111111111111111011","000000000000000101","111111111111101001","000000000000010110","111111111111110110","000000000000010011","111111111111111101","000000000000001001","000000000000000000","000000000000101010","111111111111110011","111111111111111100","111111111111011011","000000000000011110","000000000000101010","111111111111100001","111111111111110110","000000000000000111","111111111111100001","111111111111100101","111111111111101011","111111111111100000","111111111111100010","000000000000101011","111111111111011110","000000000000001001","000000000000001110","000000000000010111","000000000000011100","000000000000010000","000000000000111001","111111111111110010","111111111111110011","000000000000011100","000000000000000010","000000000000000001","000000000000010001","000000000000001001","000000000000001001","111111111111111011","111111111111100110","111111111111100100","000000000000101110","111111111111110110","111111111111111111","111111111111111000","000000000000010100","000000000000010110","000000000000001111","000000000000100001","111111111111011101","000000000000010011","000000000000010111","111111111111011111","111111111111110101","000000000000001011","111111111111001101","111111111111111000","000000000000010011","111111111111111100","111111111111110100","111111111111110100","111111111111010101","111111111111011101","111111111111111110","000000000000101011","000000000000101111","111111111111110110","000000000000100011","000000000000011000","000000000000001110","111111111111111100","000000000000010000","000000000000011111","111111111111111010","000000000000010101","111111111111001100","111111111111111011","111111111111100100","000000000000101001","000000000000001110","111111111111110011","000000000000101001","111111111111010000","000000000000011111","000000000000100111","000000000000000001","000000000000101001","000000000000010100","111111111111111111","111111111111110001","111111111111011001","111111111111101101","000000000000001000","000000000000101000","000000000000011001","111111111111110000","111111111111100011","111111111111110010","000000000000001001","000000000000010100","000000000000011010","111111111111111100","111111111111111101","111111111111110110","111111111111100100","000000000000000010","111111111111100111","111111111111101110","111111111111111110","000000000000100001","000000000000101001","000000000000001000","000000000000000010","000000000000110101","000000000000000010","111111111111111011","000000000000011111","000000000000011110","000000000000001100","111111111111010001","111111111111111001","111111111111001010","111111111111110000","000000000000010001","111111111111111100"),
("000000000000001100","111111111110111011","111111111111101110","000000000000000111","111111111111100010","000000000000010101","111111111111011111","000000000000001100","000000000000011110","111111111111100101","000000000000000101","000000000000000111","111111111111110100","111111111111100111","111111111111100100","000000000000010010","000000000000001101","000000000000000111","000000000000011110","000000000000010000","000000000000010100","111111111111111111","111111111111010101","111111111111011000","111111111111111100","000000000000010000","111111111111110110","111111111111110110","111111111111110100","000000000000010010","000000000000100111","000000000000011110","111111111111111110","111111111111111010","000000000000011111","111111111111110000","000000000000001000","000000000000100000","000000000000000101","000000000000001110","000000000000001110","000000000000001110","111111111111110110","111111111111001001","000000000000000000","111111111111110101","111111111111101011","111111111111101110","000000000000010011","000000000000010101","000000000000000010","000000000000000101","000000000000010111","000000000000011111","111111111111111111","111111111111101011","111111111111100001","111111111111111110","111111111111010101","000000000000010001","000000000000001011","111111111111111010","111111111111010110","111111111111100000","111111111111000100","000000000000000000","000000000000001001","000000000000010000","000000000000110000","111111111111110001","111111111111111100","000000000000011110","111111111111101100","000000000000000110","000000000000000110","000000000000011101","000000000000001011","111111111111111010","111111111111100110","000000000000000111","111111111111010110","000000000000001100","111111111111011101","000000000000011001","000000000000001011","111111111111101111","000000000000101010","000000000000101101","000000000000001111","000000000000011110","000000000000000011","111111111111011111","111111111111111101","111111111111001010","000000000000000111","111111111111110000","000000000000011001","000000000000001011","111111111111011101","111111111111111010","111111111111110110","000000000000000110","111111111111100111","111111111111111010","111111111111101100","000000000000001000","000000000000000000","111111111111110101","000000000000001111","111111111111100001","111111111111110000","111111111111101000","000000000000010000","000000000000000011","000000000000100010","111111111111101000","000000000000000011","000000000000000001","000000000000000110","000000000000000100","000000000000011010","000000000000000001","111111111111100111","000000000000001110","111111111111010010","111111111111110111","000000000000000111","000000000000000001"),
("111111111111111111","111111111111001000","111111111111110100","000000000000000110","111111111111101001","111111111111110110","111111111111101101","111111111111111010","000000000000000010","111111111111111110","111111111111110010","000000000000001001","000000000000001010","000000000000010101","111111111111011001","111111111111110011","000000000000000001","000000000000010101","000000000000001110","111111111111111101","000000000000001000","000000000000111000","000000000000000000","111111111111011010","111111111111110000","111111111111111111","111111111111011011","111111111111110110","000000000000001100","000000000000001001","000000000000010100","000000000000011010","000000000000001010","111111111111101101","000000000000010101","000000000000000010","000000000000010010","000000000000010101","000000000000100001","000000000000001000","000000000000001110","000000000000101010","000000000000000101","111111111111011011","111111111111101010","111111111111110000","111111111111011001","000000000000000111","000000000000010110","000000000000001100","000000000000001010","000000000000001011","111111111111111011","000000000000000010","000000000000001110","111111111111101010","111111111111101011","000000000000010010","111111111111101100","000000000000010010","000000000000010010","000000000000011010","111111111111100101","111111111111100011","111111111111001011","000000000000000000","111111111111101110","000000000000100110","000000000000010011","000000000000000101","000000000000000000","000000000000011010","111111111111110100","111111111111111100","000000000000001100","000000000000011000","000000000000010000","111111111111101111","111111111111111111","111111111111110111","000000000000000000","111111111111110110","000000000000000000","000000000000011001","000000000000001001","111111111111100010","000000000000001010","000000000000011010","111111111111110000","111111111111110001","111111111111111110","111111111111111110","111111111111010010","111111111111011100","111111111111111000","000000000000001101","111111111111100001","111111111111110110","111111111111100111","111111111111111010","111111111111100111","111111111111110101","111111111111101111","111111111111111010","111111111111111001","111111111111110100","111111111111101100","000000000000001101","000000000000011011","111111111111100001","111111111111110000","111111111111111001","111111111111111001","000000000000001000","111111111111101000","111111111111111001","111111111111110000","000000000000000000","000000000000000111","000000000000001110","000000000000101011","111111111111111011","111111111111011000","111111111111100010","111111111111101110","111111111111100110","000000000000000100","111111111111111010"),
("111111111111101111","111111111111100100","111111111111111101","111111111111111110","111111111111111010","111111111111111011","000000000000001010","111111111111111101","111111111111110110","111111111111110111","000000000000010101","111111111111111110","000000000000001101","000000000000101001","111111111111001101","000000000000010001","000000000000000110","111111111111111111","000000000000000100","000000000000101011","000000000000000000","000000000000101110","000000000000101001","000000000000001000","111111111111100110","111111111111100011","111111111111111001","111111111111110000","111111111111111110","000000000000010001","111111111111100000","000000000000010100","111111111111111000","111111111111011100","000000000000010011","000000000000001010","000000000000000001","000000000000001001","000000000000011111","111111111111110010","111111111111110011","111111111111111101","111111111111100001","111111111110110101","111111111111100100","111111111111111100","000000000000000010","111111111111101011","000000000000000000","111111111111111101","000000000000011011","000000000000001100","000000000000000001","000000000000010011","000000000000000000","111111111111110101","111111111111011111","000000000000100100","111111111111111011","000000000000000110","000000000000001100","000000000000010010","000000000000000100","111111111111110001","111111111110101010","111111111111101101","000000000000000111","000000000000001001","000000000000111001","000000000000010000","000000000000000010","000000000000010111","111111111111011001","111111111111110011","111111111111101110","000000000000110101","000000000000001000","000000000000001101","000000000000001001","000000000000000000","111111111111111110","111111111111101101","000000000000000111","000000000000001011","000000000000011000","111111111111110101","000000000000001110","000000000000000010","111111111111111000","111111111111111111","000000000000000010","000000000000000100","111111111111011111","111111111111110110","111111111111100110","000000000000100000","111111111111010110","000000000000000001","111111111111001100","111111111111111010","111111111111011101","111111111111111010","111111111111110000","111111111111111001","111111111111111000","000000000000001101","111111111111101110","000000000000000111","000000000000011100","000000000000000000","000000000000000110","000000000000000010","111111111111011101","000000000000000100","000000000000001100","000000000000001100","111111111111101010","000000000000001010","000000000000000111","000000000000011101","000000000000101000","111111111111111100","111111111111010101","000000000000001101","111111111111101111","111111111111111001","000000000000010100","111111111111110001"),
("111111111111101110","111111111111011011","111111111111101111","000000000000010011","111111111111101011","111111111111101000","000000000000000111","000000000000000000","000000000000011111","111111111111111101","000000000000001010","111111111111111100","000000000000011110","000000000000010000","111111111111011110","000000000000001001","000000000000010001","000000000000000111","111111111111111011","000000000000000111","000000000000000110","000000000001000100","000000000000001011","000000000000001001","111111111111111111","111111111111111011","111111111111101011","111111111111111100","000000000000010110","000000000000000000","111111111111100110","000000000000000101","111111111111111001","111111111111011111","111111111111101001","000000000000000010","000000000000001000","111111111111111100","000000000000101111","111111111111111111","000000000000000110","111111111111111000","111111111111011001","111111111111011001","111111111111101011","000000000000001011","111111111111011011","111111111111011010","000000000000001101","111111111111111001","000000000000010000","111111111111111101","111111111111111110","000000000000001110","111111111111111111","000000000000010101","111111111111100011","000000000000001000","000000000000101011","111111111111101111","000000000000000001","000000000000000001","000000000000010111","000000000000010001","111111111111011011","000000000000001101","000000000000001101","000000000000000100","000000000000100000","000000000000000011","000000000000001100","000000000000010100","111111111110111101","111111111111101101","111111111111110010","000000000000100001","111111111111101101","000000000000011100","000000000000011011","000000000000001110","111111111111110101","000000000000000000","000000000000100010","000000000000001001","000000000000011100","000000000000100100","000000000000011011","111111111111101110","111111111111110100","000000000000011001","000000000000001000","111111111111111011","111111111111101001","111111111111110000","111111111111011100","000000000000010100","000000000000001010","111111111111111011","111111111111100101","000000000000011010","111111111111011110","111111111111101101","000000000000000111","000000000000010011","111111111111111000","111111111111111110","111111111111110001","111111111111110001","000000000000101000","000000000000001110","000000000000001011","000000000000010100","111111111111100011","111111111111111001","111111111111111101","000000000000001000","111111111111101100","000000000000001110","000000000000000101","000000000000100010","000000000000000001","111111111111110101","111111111111111101","000000000000000101","111111111111111101","111111111111010100","000000000000010010","000000000000000100"),
("111111111111111000","111111111110111100","111111111111110011","000000000000001101","111111111111110001","111111111111110110","000000000000100111","000000000000001100","111111111111111111","111111111111111001","000000000000001000","111111111111111000","111111111111111001","111111111111111110","111111111111010000","000000000000010010","000000000000001101","000000000000010100","000000000000001001","000000000000000111","000000000000000011","000000000001000100","111111111111111110","000000000000010111","111111111111110110","000000000000011011","000000000000001111","111111111111111011","000000000000001001","000000000000001001","111111111111101110","111111111111111001","000000000000001010","111111111111010111","111111111111100100","000000000000010011","000000000000000000","111111111111101011","000000000000011101","111111111111101010","000000000000000010","000000000000000111","111111111111010100","111111111111101010","000000000000000011","111111111111110110","111111111111100111","000000000000001011","111111111111111010","111111111111110011","000000000000010011","000000000000100101","111111111111111011","111111111111111101","111111111111111110","000000000000000000","111111111111011010","111111111111111011","000000000000000010","000000000000000000","111111111111011101","111111111111100101","000000000000001000","000000000000000100","000000000000010000","000000000000010010","000000000000010111","111111111111111011","111111111111111100","111111111111111101","111111111111110111","111111111111111101","111111111111101000","111111111111011110","111111111111101101","000000000000110111","000000000000001000","000000000000100000","111111111111110100","000000000000011110","111111111111111111","000000000000011101","000000000000000000","111111111111110010","000000000000001101","000000000000001000","000000000000000010","000000000000000100","111111111111110110","000000000000001001","111111111111101111","000000000000100101","000000000000011000","111111111111110001","111111111111011011","000000000000010100","000000000000010101","000000000000010100","111111111111100110","000000000000000111","111111111111011010","111111111111101101","000000000000000101","000000000000010001","000000000000001000","000000000000011011","000000000000010110","000000000000000000","000000000000011011","111111111111110110","000000000000010001","000000000000010111","111111111111111011","111111111111110010","111111111111110111","000000000000000110","000000000000001111","000000000000001000","000000000000010110","000000000000010001","000000000000000001","000000000000011000","111111111111110100","000000000000011101","111111111111110110","111111111111011110","111111111111111111","111111111111111000"),
("111111111111011100","111111111110100001","111111111111101111","000000000000000100","000000000000011001","111111111111110101","000000000000010000","111111111111110101","000000000000000011","000000000000000011","000000000000010111","111111111111110100","111111111111110100","000000000000000100","111111111111011001","000000000000100001","111111111111101010","000000000000010011","000000000000000001","000000000000010110","000000000000010100","000000000000011111","000000000000000111","000000000000010111","000000000000000001","111111111111110010","000000000000011011","000000000000011000","111111111111111100","000000000000100100","111111111111111000","111111111111101000","000000000000010101","111111111111011101","111111111111110100","000000000000000000","111111111111110101","000000000000001110","000000000000010110","111111111111111001","000000000000001101","000000000000011001","111111111111100110","000000000000000001","000000000000001111","000000000000000110","111111111111111011","111111111111111000","000000000000000000","111111111111100101","000000000000100110","000000000000000101","000000000000000000","111111111111110010","000000000000001001","000000000000000110","111111111111101100","000000000000010111","000000000000001011","111111111111110110","111111111111101000","111111111111110000","111111111111111011","000000000000010000","111111111111111110","111111111111111101","000000000000100000","000000000000001110","000000000000001001","000000000000011000","111111111111110011","000000000000001111","111111111111101010","000000000000000101","111111111111101110","000000000000011111","000000000000001110","000000000000010101","111111111111101100","000000000000000000","000000000000000100","000000000000000111","111111111111011001","000000000000000000","000000000000010000","000000000000000000","111111111111111111","000000000000000101","111111111111110101","000000000000010011","000000000000000001","000000000000001011","000000000000000010","000000000000000110","111111111111010110","000000000000001001","000000000000011011","000000000000000000","000000000000000101","111111111111101000","111111111111100010","111111111111100100","000000000000001110","000000000000100111","000000000000001101","000000000000001101","000000000000000001","111111111111110111","000000000000010101","000000000000010110","000000000000000010","000000000000000010","111111111111110110","111111111111101000","111111111111111000","000000000000010010","000000000000000000","000000000000100101","111111111111110111","111111111111111000","111111111111111100","000000000000010001","000000000000001110","000000000000001010","111111111111110100","111111111111100100","000000000000000010","111111111111011010"),
("111111111111111100","111111111111010010","000000000000011100","000000000000001111","000000000000001000","111111111111110001","000000000000011111","000000000000000110","000000000000001000","000000000000010000","000000000000001110","111111111111111100","111111111111110010","000000000000010010","111111111111110101","000000000000001011","000000000000000000","000000000000001010","000000000000000000","000000000000000101","111111111111110101","111111111111111110","000000000000011100","000000000000001011","000000000000011101","000000000000000001","000000000000100000","000000000000011001","111111111111101101","000000000000110010","111111111111111010","111111111111110011","000000000000001101","000000000000000000","000000000000000001","000000000000010000","111111111111111100","000000000000001011","000000000000001100","000000000000011100","000000000000011011","111111111111110110","111111111111100001","111111111111111001","111111111111111111","000000000000000011","000000000000000011","111111111111101100","000000000000010111","111111111111101011","000000000000000011","000000000000010101","111111111111111101","000000000000011001","000000000000001001","111111111111110110","111111111111110101","111111111111111110","000000000000010010","111111111111101111","111111111111111110","111111111111111001","000000000000100000","000000000000000111","000000000000011010","000000000000000000","000000000000010000","111111111111111110","000000000000000100","000000000000001011","111111111111111101","111111111111111010","111111111111110000","000000000000001001","111111111111111010","000000000000111010","111111111111110110","111111111111111001","000000000000000111","000000000000100010","000000000000000110","111111111111111100","111111111111001101","000000000000000110","000000000000010110","000000000000000000","000000000000011110","000000000000010110","000000000000000010","000000000000001000","111111111111101011","000000000000011000","000000000000000010","000000000000001010","111111111111011101","000000000000101010","000000000000100000","111111111111101100","000000000000011010","000000000000010001","111111111111111001","000000000000000000","111111111111111111","000000000000000110","000000000000000111","000000000000000001","111111111111110100","111111111111100011","000000000000001011","000000000000001010","000000000000001010","000000000000100101","000000000000010101","111111111111111110","111111111111101101","000000000000011011","111111111111111100","000000000000011001","000000000000100101","000000000000100101","000000000000001000","000000000000001011","000000000000001011","111111111111110001","111111111111111011","111111111111100111","000000000000100001","111111111111111111"),
("111111111111110101","111111111111001110","000000000000000101","000000000000001010","111111111111111101","111111111111100111","000000000000000100","111111111111110111","000000000000001111","000000000000000011","000000000000011010","111111111111110101","111111111111101000","111111111111101000","111111111111111100","000000000000101100","111111111111110100","000000000000001011","000000000000000101","000000000000010000","000000000000001000","111111111111101001","000000000000001111","000000000000001011","000000000000001110","111111111111101000","000000000000010000","000000000000100001","111111111111110000","000000000000010101","111111111111110110","111111111111110010","000000000000001011","111111111111110010","111111111111101011","000000000000010000","111111111111110101","111111111111111101","000000000000000000","111111111111111001","000000000000001101","111111111111111100","000000000000000101","111111111111111100","000000000000011110","000000000000000010","000000000000011100","111111111111010001","111111111111111011","000000000000000000","111111111111111000","000000000000110000","000000000000010011","000000000000010111","000000000000000100","000000000000001011","000000000000000000","000000000000000110","000000000000010010","000000000000010001","000000000000000101","000000000000000010","000000000000100111","000000000000011000","000000000000001100","000000000000001010","000000000000001011","000000000000010111","111111111111110111","000000000000000001","111111111111111010","000000000000010010","111111111111101110","000000000000010011","111111111111100101","000000000000011110","000000000000000110","000000000000001001","000000000000000101","000000000000011001","111111111111110100","000000000000000000","111111111111101100","000000000000010010","000000000000100100","111111111111110101","000000000000011100","000000000000000100","111111111111110110","000000000000010000","111111111111110111","000000000000000101","111111111111100011","000000000000000001","111111111111100111","000000000000000100","000000000000001111","000000000000001011","000000000000010100","000000000000011001","000000000000000001","111111111111110100","000000000000100110","000000000000011101","000000000000010010","000000000000010110","000000000000001001","111111111111110101","111111111111101111","111111111111110111","111111111111110010","000000000000010100","000000000000010000","111111111111111011","111111111111101001","111111111111111100","000000000000000100","000000000000101111","000000000000100110","000000000000110000","000000000000010100","000000000000011110","111111111111110010","111111111111101010","000000000000010010","111111111111101001","000000000000000101","000000000000010111"),
("111111111111111110","111111111111011111","111111111111111001","000000000000001101","000000000000000101","111111111111110000","000000000000100101","111111111111100110","111111111111101110","000000000000000101","000000000000101000","000000000000000101","111111111111110101","111111111111101100","111111111111110010","000000000000011001","000000000000010010","000000000000010011","000000000000001001","000000000000001010","000000000000010011","111111111111010101","111111111111111111","000000000000110101","000000000000010100","000000000000010001","000000000000001110","000000000000011010","111111111111110001","000000000000110011","000000000000000011","111111111111110001","000000000000000000","000000000000010110","111111111111110001","111111111111111011","111111111111101010","111111111111101011","111111111111110110","111111111111110000","000000000000000111","000000000000011111","000000000000000111","000000000000011010","000000000000001010","000000000000010000","000000000000001010","111111111111111000","000000000000000010","111111111111111001","111111111111111111","000000000000000110","000000000000001010","000000000000001000","000000000000000101","000000000000001001","111111111111110011","000000000000001000","000000000000001000","111111111111111000","111111111111110111","111111111111110010","000000000000001011","000000000000000010","000000000000000111","111111111111111011","000000000000000000","000000000000001110","000000000000000101","000000000000000000","000000000000000101","111111111111110011","111111111111100111","111111111111110110","111111111111100011","000000000000010111","000000000000001111","111111111111111011","111111111111111011","000000000000010000","000000000000011010","000000000000000000","111111111111101100","000000000000001110","000000000000100101","111111111111101111","000000000000011001","000000000000001001","111111111111110011","000000000000001100","111111111111101011","000000000000011110","111111111111111011","000000000000011011","111111111111101111","000000000000000101","000000000000011100","111111111111011110","111111111111111101","111111111111111101","111111111111111110","000000000000010001","000000000000100100","000000000000001000","000000000000001010","000000000000010000","000000000000010011","111111111111101111","111111111111011010","111111111111110010","000000000000000110","000000000000110011","111111111111111111","000000000000001010","111111111111011011","111111111111111110","000000000000000100","000000000000001100","000000000000001101","000000000000010010","000000000000000001","000000000000010110","000000000000001111","000000000000001001","111111111111101011","111111111111111001","000000000000001101","111111111111111000"),
("111111111111101101","111111111111110110","111111111111111111","000000000000010000","000000000000001101","111111111111101100","000000000000001100","111111111111100100","111111111111110111","000000000000010001","000000000000011011","000000000000010110","000000000000000001","111111111111100110","111111111111101110","000000000000010000","000000000000001001","000000000000001101","000000000000010011","111111111111111100","000000000000011111","111111111111100010","000000000000000111","000000000000001001","000000000000000000","111111111111110001","000000000000011101","000000000000010010","000000000000001110","000000000000011100","111111111111100110","111111111111011010","111111111111111111","000000000000011011","000000000000000100","000000000000000000","111111111111111111","111111111111111100","111111111111110100","111111111111111010","111111111111111101","111111111111111110","000000000000010001","000000000000011010","000000000000000110","111111111111111010","000000000000011010","111111111111011101","000000000000000111","111111111111110111","111111111111100011","000000000000100110","000000000000000101","111111111111110000","111111111111110011","111111111111101011","000000000000010100","000000000000011011","111111111111110100","111111111111111001","111111111111111111","000000000000010101","000000000000000011","000000000000010110","111111111111111011","000000000000010001","111111111111110100","111111111111111110","111111111111101111","000000000000001011","000000000000000000","111111111111110101","111111111111011110","111111111111111100","000000000000000000","000000000000000101","000000000000001001","111111111111111000","000000000000000010","111111111111111111","111111111111111001","111111111111111101","111111111111101101","000000000000010011","000000000000010101","111111111111011101","000000000000010100","111111111111100101","000000000000001001","000000000000000100","000000000000000001","000000000000101000","111111111111110010","000000000000000111","000000000000000000","111111111111110100","000000000000000000","111111111111111011","111111111111110100","111111111111101010","111111111111110001","000000000000011100","000000000000010110","000000000000011011","000000000000011001","000000000000011101","111111111111111110","111111111111110010","111111111111111101","000000000000000100","000000000000010110","000000000000001000","000000000000001100","000000000000011011","000000000000010011","000000000000001000","000000000000000001","000000000000000010","000000000000011110","000000000000001110","000000000000001101","111111111111110001","111111111111111111","111111111111101100","111111111111101011","000000000000000000","000000000000011011","000000000000001000"),
("000000000000010000","000000000000010000","000000000000010001","000000000000001110","000000000000001100","000000000000000011","111111111111110101","111111111111011100","111111111111110111","000000000000001111","000000000000001011","000000000000110011","000000000000000101","111111111111100101","000000000000001101","000000000000001010","111111111111110011","111111111111111011","000000000000000100","111111111111110101","000000000000000000","111111111111011000","000000000000000000","000000000000000010","000000000000000101","111111111111110001","000000000000010101","000000000000000100","111111111111111101","000000000000100110","111111111111101101","111111111111111100","000000000000001100","000000000000010101","111111111111110010","000000000000000010","111111111111111100","000000000000000000","111111111111110110","111111111111111101","111111111111111000","000000000000001100","000000000000010010","000000000000000101","000000000000011110","000000000000001001","000000000000001100","111111111111100111","000000000000010110","111111111111111000","111111111111100110","000000000000001110","000000000000000101","111111111111110000","000000000000001101","111111111111110010","000000000000010101","000000000000001011","111111111111111110","111111111111101110","111111111111110000","000000000000001000","111111111111101110","000000000000010101","111111111111101110","000000000000011000","111111111111110000","111111111111111000","111111111111110111","000000000000010111","111111111111110000","000000000000010001","111111111111101000","000000000000000101","111111111111111001","000000000000000011","111111111111101101","111111111111111101","111111111111110100","000000000000010100","111111111111111101","000000000000011001","111111111111101010","111111111111111100","000000000000010110","111111111111111111","000000000000011010","111111111111101010","000000000000000111","111111111111101100","000000000000010110","000000000000100011","000000000000000001","111111111111111110","000000000000000010","111111111111101000","111111111111111110","000000000000000111","111111111111110100","111111111111100110","111111111111011111","000000000000010101","000000000000011010","000000000000010010","111111111111111100","000000000000000001","000000000000010010","111111111111110111","111111111111111010","111111111111111000","000000000000001000","000000000000100100","000000000000011010","000000000000001100","000000000000001111","000000000000000000","000000000000001111","000000000000001111","000000000000001010","000000000000011110","000000000000001100","111111111111110110","000000000000001100","000000000000000000","111111111111100001","000000000000011000","000000000000011000","000000000000010110"),
("000000000000000110","000000000000101000","111111111111101010","000000000000000011","000000000000011110","111111111111110100","111111111111011010","111111111111111110","111111111111110010","111111111111111110","000000000000000110","000000000000111010","111111111111110111","111111111111110100","000000000000000000","000000000000000110","111111111111101001","111111111111111100","000000000000010001","111111111111110010","000000000000100000","000000000000001101","000000000000000000","000000000000010000","111111111111111110","000000000000000101","000000000000011111","111111111111111011","000000000000001111","000000000000100010","111111111111100011","111111111111111100","000000000000001011","000000000000001101","111111111111110010","000000000000010010","111111111111101010","111111111111111100","111111111111110110","000000000000001111","000000000000011000","000000000000011000","000000000000100000","000000000000011001","000000000000000001","111111111111011010","000000000000001100","111111111111110101","000000000000001101","000000000000001100","111111111111111011","111111111111111100","000000000000001111","111111111111110110","111111111111110010","111111111111101100","000000000000001010","000000000000001000","111111111111111100","000000000000000010","000000000000001011","111111111111110011","111111111111101110","111111111111111101","000000000000000111","000000000000000111","111111111111010100","111111111111111111","111111111111111100","000000000000001011","000000000000000011","000000000000010111","111111111111110001","111111111111111010","111111111111110001","111111111111110010","111111111111110010","000000000000010100","000000000000000111","000000000000000011","000000000000011101","000000000000010110","111111111111011111","111111111111101101","000000000000101010","111111111111110010","000000000000011110","000000000000000011","000000000000001010","111111111111110111","000000000000011010","000000000000011011","000000000000000111","000000000000000111","000000000000001100","111111111111111110","111111111111111001","111111111111110000","000000000000000111","111111111111110001","111111111111110010","000000000000010101","111111111111110011","000000000000011100","111111111111111011","111111111111110000","111111111111111100","111111111111110111","000000000000001100","111111111111110010","000000000000000000","000000000000010001","000000000000001101","000000000000011110","000000000000000100","000000000000001010","111111111111111111","000000000000001110","111111111111110011","111111111111111111","000000000000001111","000000000000000110","000000000000000000","000000000000010001","111111111111011101","000000000000010110","000000000000001110","111111111111111010"),
("000000000000011001","000000000000011001","000000000000000110","000000000000011001","000000000000000100","000000000000000000","111111111111110101","111111111111111100","111111111111111110","111111111111111011","000000000000110000","000000000000101001","000000000000000000","111111111111100010","111111111111111001","000000000000011101","111111111111101010","000000000000000110","111111111111111010","000000000000001100","000000000000010110","000000000000001101","000000000000010100","111111111111111100","000000000000000010","000000000000001001","000000000000011001","000000000000010011","000000000000001010","111111111111111011","111111111111111000","111111111111101100","111111111111110011","000000000000000100","111111111111110111","000000000000010101","111111111111110000","000000000000000011","000000000000011111","000000000000001111","111111111111111000","000000000000010001","111111111111111001","000000000000001000","000000000000001101","111111111111100111","000000000000100000","111111111111100011","000000000000010111","111111111111111101","111111111111101000","000000000000010001","111111111111111010","000000000000001000","111111111111110000","000000000000000001","000000000000001010","111111111111110010","111111111111110100","111111111111110011","111111111111100001","111111111111110110","111111111111101000","111111111111111011","111111111111111000","000000000000001110","111111111110110100","000000000000000011","111111111111110000","111111111111111110","111111111111111100","000000000000001100","111111111111101011","000000000000000101","111111111111111110","111111111111110100","000000000000010001","000000000000001100","111111111111100110","111111111111111011","000000000000000100","000000000000001001","111111111111010111","111111111111111011","000000000000100001","111111111111101100","000000000000011000","000000000000001000","000000000000010110","111111111111101100","000000000000010111","000000000000010111","000000000000001110","111111111111111101","000000000000000111","111111111111101001","000000000000000101","000000000000001001","111111111111010100","111111111111101100","111111111111010100","000000000000100001","111111111111100100","000000000000001101","000000000000000011","000000000000010011","111111111111111111","111111111111110000","000000000000000011","111111111111110100","111111111111111001","000000000000001010","000000000000001111","111111111111111011","000000000000001000","000000000000000011","111111111111111111","000000000000000001","000000000000000110","000000000000000010","000000000000000011","111111111111111001","111111111111111111","000000000000001001","111111111111110100","000000000000001100","000000000000011001","000000000000001000"),
("000000000000010000","000000000000101010","111111111111110011","000000000000000101","000000000000010111","000000000000001011","111111111111101001","000000000000011100","111111111111110111","111111111111111100","000000000000011100","000000000000110011","111111111111110100","111111111111010100","000000000000001011","000000000000001101","111111111111100110","111111111111110110","111111111111111001","111111111111110111","000000000000010111","000000000000100000","111111111111110110","111111111111011010","000000000000001011","000000000000000100","000000000000011011","111111111111110101","111111111111111111","000000000000001110","000000000000010001","111111111111110101","111111111111110011","000000000000001000","111111111111100110","000000000000010100","111111111111100110","111111111111111100","000000000000010011","111111111111110000","000000000000011001","111111111111101111","000000000000000000","000000000000101000","000000000000011110","000000000000000010","111111111111110011","111111111111100101","111111111111110111","111111111111111011","111111111111100000","000000000000001001","111111111111100100","000000000000000000","111111111111101101","000000000000001110","111111111111111001","000000000000000101","111111111111111111","111111111111111000","111111111111101101","000000000000000001","111111111111100011","000000000000001010","000000000000110000","111111111111111111","111111111110110100","111111111111111000","111111111111101011","000000000000000001","000000000000010011","000000000000011101","111111111111100001","000000000000001101","000000000000000101","111111111111100000","111111111111101110","000000000000011101","111111111111111101","111111111111101001","000000000000000110","000000000000000101","111111111111001010","111111111111100011","000000000000010001","111111111111101010","000000000000010110","111111111111101110","000000000000000010","111111111111101100","000000000000001111","000000000000001011","111111111111111011","000000000000000000","000000000000001111","111111111111001101","111111111111111000","000000000000000001","111111111111010100","111111111111101101","111111111111101001","111111111111111000","111111111111110111","000000000000011111","111111111111101100","000000000000011000","000000000000000010","111111111111111011","111111111111110111","000000000000001010","000000000000010000","000000000000001011","000000000000001101","000000000000010100","000000000000010110","111111111111101100","000000000000000100","000000000000000000","000000000000001111","000000000000001111","000000000000001111","111111111111111000","111111111111110000","000000000000100110","111111111111010000","000000000000010110","000000000000000100","000000000000011101"),
("111111111111111111","000000000000101011","111111111111100111","000000000000000000","000000000000100111","000000000000100000","111111111111101001","000000000000011000","111111111111110111","000000000000000001","000000000000011100","000000000000100000","111111111111110011","111111111111011100","111111111111110011","000000000000010011","000000000000000100","000000000000000110","111111111111111111","111111111111110000","111111111111111000","000000000000011101","000000000000010000","111111111111101001","111111111111110010","000000000000111100","111111111111110110","111111111111111100","111111111111110000","111111111111111110","111111111111110101","111111111111011110","000000000000000010","111111111111111010","000000000000001011","000000000000011101","111111111111110001","000000000000001001","000000000000001101","000000000000010100","111111111111111100","111111111111101111","000000000000001111","000000000000100001","000000000000111001","111111111111111000","111111111111111000","111111111111100011","000000000000001101","000000000000001001","111111111111101111","000000000000001000","111111111111100001","000000000000001110","111111111111101011","000000000000000101","111111111111101010","111111111111111010","111111111111101001","000000000000000010","111111111111011111","000000000000001111","111111111111011110","000000000000001101","000000000000100011","111111111111100101","111111111110100101","000000000000100000","111111111111101000","111111111111101011","000000000000011000","000000000000000111","111111111111100111","111111111111111111","000000000000101100","111111111111101001","111111111111111101","000000000000010011","000000000000000000","000000000000000000","000000000000000111","000000000000011000","111111111111011110","111111111111100110","000000000000000101","111111111111101100","000000000000000001","000000000000000011","000000000000110110","111111111111111010","111111111111110101","000000000000000111","111111111111100101","111111111111101000","111111111111111100","111111111111101110","111111111111111100","000000000000101001","111111111111010100","111111111111101011","000000000000000010","111111111111110101","111111111111010001","000000000000000110","111111111111100111","000000000000001010","111111111111111111","111111111111010110","000000000000000000","111111111111111111","000000000000000000","000000000000010000","000000000000110010","000000000000001011","111111111111110110","111111111111101110","000000000000001100","111111111111111100","111111111111100010","111111111111111100","000000000000000100","111111111111111110","111111111111111101","000000000000011110","111111111110111000","000000000000010100","111111111111111110","000000000000100001"),
("000000000000010001","000000000000010000","000000000000001001","000000000000000000","000000000000100001","000000000000110000","111111111111100100","000000000000011100","000000000000000011","000000000000010000","000000000000110100","111111111111111010","111111111111111001","111111111111100001","000000000000000010","000000000000010011","000000000000000010","111111111111110001","000000000000001001","000000000000000011","111111111111011110","000000000000011100","000000000000001101","111111111111001100","111111111111111000","000000000000100111","000000000000001111","000000000000010110","111111111111111011","111111111111101001","000000000000011000","111111111111111001","111111111111100100","111111111111111100","000000000000001010","000000000000000111","111111111111100110","000000000000000010","000000000000001010","000000000000000000","111111111111111000","111111111111011111","000000000000001100","000000000000010010","000000000000101100","111111111111111000","000000000000001101","000000000000000011","111111111111110000","111111111111100100","000000000000000001","111111111111111100","111111111111100110","000000000000001010","111111111111111111","000000000000010000","111111111111011001","000000000000000011","111111111111100000","000000000000010001","111111111111010001","111111111111110010","000000000000000011","000000000000001010","111111111111110101","111111111111101100","111111111110110001","000000000000000101","111111111111011111","111111111111110101","000000000000011010","000000000000000000","111111111110111000","111111111111100101","000000000000101000","111111111111100010","000000000000100001","000000000000000011","000000000000000011","111111111111111011","000000000000010010","000000000000001100","111111111111010010","111111111110111101","111111111111111101","111111111111110000","000000000000001000","000000000000000101","000000000000010100","111111111111111000","111111111111111110","000000000000000011","111111111111101101","111111111111101110","111111111111110101","111111111111100100","111111111111111010","000000000000010001","111111111111110010","111111111111100000","111111111111111110","000000000000000010","111111111111011011","000000000000000000","111111111111111101","111111111111111010","111111111111111010","111111111111011101","000000000000011110","111111111111111100","000000000000010110","000000000000000101","000000000000001100","000000000000000000","111111111111100100","111111111111110011","111111111111110100","111111111111111100","111111111111101011","111111111111110001","111111111111111010","000000000000000010","111111111111111000","000000000000100110","111111111111001100","000000000000001000","000000000000001111","000000000000001001"),
("111111111111111101","000000000000010101","000000000000000111","000000000000000111","000000000000011110","000000000000011011","111111111111111000","000000000000011000","000000000000000100","000000000000010010","000000000000011100","111111111111110000","111111111111110101","111111111111101011","000000000000000001","000000000000000010","111111111111110011","000000000000000000","000000000000000110","111111111111111011","111111111111101010","000000000000001010","111111111111110100","111111111111010011","111111111111101110","000000000000010100","111111111111110001","000000000000011101","111111111111110000","111111111111111010","000000000000001000","111111111111100100","000000000000001010","111111111111101110","000000000000001001","000000000000001100","111111111111101010","000000000000000000","111111111111110110","111111111111100101","000000000000000010","111111111111101000","000000000000000000","000000000000101101","000000000000010100","111111111111100101","000000000000000101","000000000000000100","111111111111110000","111111111111110100","111111111111011000","000000000000001010","111111111111100100","000000000000011100","111111111111101101","000000000000010010","111111111111001101","000000000000000000","111111111111011101","000000000000010011","111111111111001111","000000000000000000","111111111111101000","000000000000000000","111111111111010110","111111111111111011","111111111111010000","111111111111110101","111111111111101100","111111111111101010","000000000000100010","000000000000000101","111111111111100011","111111111111011110","000000000000110001","111111111111100001","000000000000000111","000000000000011100","000000000000001011","111111111111101111","000000000000001000","000000000000011101","111111111111110000","111111111111110010","111111111111111101","000000000000000100","111111111111111010","000000000000000100","111111111111110100","111111111111101100","111111111111110010","111111111111100001","000000000000000001","111111111111010110","111111111111110001","111111111111011111","111111111111111100","111111111111111111","111111111111101000","111111111111110000","000000000000001010","111111111111111100","111111111111010111","000000000000010010","111111111111110001","111111111111111111","000000000000010111","111111111111110011","111111111111101010","111111111111011000","000000000000000110","000000000000011000","000000000000011011","111111111111110101","111111111111111000","111111111111100001","000000000000001001","111111111111100000","111111111111011110","000000000000010010","000000000000000000","111111111111111101","111111111111110000","000000000000100000","111111111111110000","000000000000000010","111111111111101111","000000000000011011"),
("000000000000000000","000000000000010101","111111111111110100","111111111111111101","000000000000100100","000000000000110010","111111111111111110","000000000000010110","000000000000011010","111111111111110111","000000000000100000","111111111111110000","000000000000010100","000000000000001111","000000000000000001","000000000000010001","000000000000001000","000000000000000011","111111111111110010","111111111111101110","111111111111001001","111111111111001100","000000000000100101","111111111111110010","111111111111110110","000000000000110000","000000000000010001","000000000000101101","111111111111100011","111111111111110011","000000000000000110","111111111111010001","000000000000001000","111111111111111101","111111111111110111","111111111111110111","111111111111111000","000000000000001110","111111111111111100","111111111111101001","111111111111111110","111111111111001010","000000000000000100","000000000000101110","000000000000100110","111111111111100100","111111111111100110","000000000000000000","111111111111101110","111111111111011000","111111111111011111","000000000000011110","111111111111011101","000000000000001110","000000000000000011","000000000000100010","111111111111100110","111111111111011100","111111111111100001","000000000000001001","111111111111010100","000000000000100010","000000000000010000","000000000000001110","111111111111110111","111111111111100111","111111111111100111","111111111111110100","111111111111010001","111111111111111111","000000000000001101","111111111111100111","111111111111010100","111111111111101100","111111111111111010","111111111111101100","000000000000010001","000000000000000000","111111111111111011","000000000000000110","000000000000000001","000000000000110000","111111111111100110","111111111111111010","111111111111101111","000000000000011101","111111111111101011","111111111111101101","000000000000000000","111111111111011101","000000000000010001","111111111111100111","111111111111110001","111111111111111110","000000000000010101","111111111111101110","000000000000000110","000000000000100010","111111111111100101","111111111111111111","111111111111111101","000000000000000001","111111111111010000","111111111111111011","111111111111100111","111111111111110101","000000000000001001","111111111111011101","111111111111011011","111111111111010111","000000000000000011","000000000000100110","000000000000000000","111111111111010101","000000000000000001","111111111111101010","111111111111111100","111111111111101001","111111111111100000","000000000000000100","000000000000001010","111111111111110010","111111111111111010","000000000000000101","111111111111110101","111111111111111100","111111111111111101","000000000000001101"),
("111111111111111011","000000000000001001","111111111111110111","000000000000100011","111111111111010001","000000000000010011","111111111111111011","000000000000110001","000000000000001001","111111111111100011","000000000000100000","111111111111110011","000000000000011000","000000000000100010","111111111111110101","000000000000011010","111111111111100000","000000000000110011","111111111111101001","000000000000000000","000000000000001111","111111111111110111","000000000000000000","111111111111100111","111111111111111100","000000000000100111","000000000000010011","000000000000100001","111111111111111110","111111111111011101","000000000000110000","111111111111111110","000000000000010101","111111111111101100","111111111111100110","111111111111111100","111111111111110011","111111111111110011","111111111111100101","111111111111010010","111111111111101000","111111111111001111","000000000000000000","000000000000001111","000000000000100000","111111111111100011","111111111111101111","000000000000001000","111111111111100000","111111111111111101","111111111111100110","000000000000100001","111111111111110001","000000000000011010","111111111111110111","000000000000010110","111111111111001111","111111111111110101","111111111111111011","000000000000000110","111111111111010000","000000000000010011","000000000000011000","000000000000000000","000000000000001010","000000000000000000","111111111111010101","111111111111101101","111111111111011100","111111111111111100","000000000000010110","111111111111101110","111111111111110011","111111111111110011","111111111111100101","111111111111111001","000000000000011001","000000000000000101","111111111111101111","111111111111110111","111111111111100000","000000000000110000","000000000000000000","111111111111101111","000000000000001110","111111111111101000","111111111111110110","111111111111111101","111111111111111011","111111111111010000","111111111111101001","000000000000000001","000000000000010000","111111111111110101","000000000000101101","111111111111101101","111111111111110100","000000000000011101","111111111111100001","000000000000000000","000000000000100110","000000000000011000","111111111111100001","000000000000010010","111111111111011110","000000000000010101","000000000000011010","111111111111110011","111111111111011001","111111111111101110","000000000000001011","000000000000001010","000000000000000100","111111111111101011","000000000000011001","111111111111110100","000000000000000000","000000000000000000","111111111111111001","111111111111111101","000000000000011000","000000000000000101","000000000000000011","000000000000001111","111111111111100010","111111111111111000","000000000000001011","000000000000000000"),
("000000000000110001","000000000000011010","000000000000010110","000000000000010010","111111111111001110","000000000000001000","111111111111111000","000000000000101110","111111111111101110","111111111111011010","000000000000101001","111111111111111011","000000000000101010","000000000000101110","111111111111111110","000000000000011010","111111111111101110","000000000000101001","111111111111100111","000000000000001110","000000000000010000","111111111111101110","111111111111100111","000000000000001000","000000000000011010","000000000000011011","000000000000000000","000000000000101001","111111111111101111","111111111111100010","000000000000111101","111111111111101010","000000000000111000","111111111111111100","111111111111111000","111111111111011001","000000000000000000","000000000000000111","111111111111100101","111111111111100000","111111111111111111","111111111111100000","000000000000000000","000000000000001010","000000000001000001","111111111111100011","111111111111100001","111111111111100001","111111111111100010","111111111111111100","111111111111011100","000000000000011010","111111111111100001","000000000000101101","000000000000001011","000000000000011000","111111111111101000","111111111111100010","111111111111110001","111111111111110010","111111111111010100","000000000000010111","000000000000000000","111111111111110100","000000000000001011","111111111111111111","111111111111100011","111111111111111101","111111111111100100","111111111111101001","000000000000001010","000000000000000001","111111111111110000","000000000000000111","000000000000000101","000000000000100101","000000000000111001","000000000000001111","111111111111101001","111111111111110010","000000000000000001","000000000000110011","111111111111110010","111111111111000111","000000000000011000","111111111111101101","000000000000000101","000000000000010100","111111111111111000","111111111111100100","111111111111101001","000000000000001010","000000000000010001","111111111111011110","000000000000010110","111111111111101101","000000000000001001","000000000000101001","000000000000000010","000000000000000001","000000000000011001","111111111111111001","000000000000001000","000000000000001001","000000000000000101","111111111111111010","000000000000001110","111111111111010001","111111111111110111","111111111111101101","000000000000001111","000000000000001001","000000000000010100","111111111111001011","000000000000001101","111111111111011000","111111111111111000","111111111111110001","111111111111110001","111111111111110111","000000000000011110","000000000000000010","000000000000010110","000000000000011010","111111111111011000","000000000000011000","000000000000010010","111111111111110110"),
("000000000000011010","000000000000010000","000000000000010100","000000000000011000","111111111111011000","111111111111101010","111111111111110111","111111111111111010","111111111111110101","111111111111100011","111111111111111111","000000000000001000","000000000000110010","000000000000100110","000000000000000011","111111111111111010","111111111111110100","000000000000010101","000000000000000111","111111111111111101","000000000000000101","000000000000010110","111111111111100010","111111111111111100","000000000000001010","000000000000000101","111111111111101111","000000000000011000","111111111111101011","000000000000001000","000000000001001111","000000000000001111","000000000000101101","000000000000000100","111111111111111011","111111111111101111","000000000000010011","000000000000010011","111111111111110101","111111111111111110","111111111111110110","111111111111110000","111111111111101000","111111111111111011","000000000000100101","111111111111100100","111111111111001101","111111111111011100","111111111111111110","111111111111101001","111111111110111001","111111111111111001","111111111111100010","000000000001000100","000000000000011101","000000000000001110","000000000000001100","000000000000001001","111111111111111011","000000000000000011","000000000000000111","000000000000001001","111111111111110110","111111111111111011","000000000000011100","000000000000000101","111111111111001000","000000000000000000","000000000000000110","000000000000000101","000000000000100000","000000000000000110","111111111111110010","111111111111111110","000000000000010011","000000000000010011","000000000000101011","000000000000011001","111111111111110110","111111111111100100","000000000000010001","000000000000101001","111111111111100001","111111111111110010","000000000000000000","000000000000001111","111111111111111010","000000000000000000","111111111111110001","000000000000001111","111111111111101110","000000000000001101","111111111111101110","111111111111000110","000000000000011001","111111111111111010","000000000000010100","000000000000111101","111111111111111101","000000000000000111","111111111111111111","111111111111100011","111111111111111110","000000000000000001","000000000000000001","111111111111011111","111111111111101111","111111111111100100","111111111111111100","111111111111100110","111111111111111111","000000000000100101","111111111111111001","111111111111111100","111111111111101011","111111111111100000","000000000000001110","111111111111011110","000000000000010001","111111111111111100","000000000000010100","000000000000001111","111111111111110010","111111111111110100","111111111111010001","000000000000001010","111111111111110010","000000000000000001"),
("000000000000001100","000000000000001001","000000000000011110","000000000000001110","111111111111111000","000000000000000001","000000000000001000","000000000000110001","000000000000001001","111111111111111101","000000000000100110","000000000000010100","111111111111110111","000000000000110010","000000000000000101","000000000000010111","111111111111011100","111111111111110100","111111111111111001","111111111111101111","111111111111110110","000000000000000011","111111111111100000","000000000000000001","111111111111111011","000000000000001000","000000000000000000","111111111111101010","000000000000000001","111111111111110100","000000000000010111","111111111111101001","000000000000000100","111111111111100101","111111111111110110","000000000000000000","000000000000000000","000000000000000011","111111111111101110","000000000000001100","111111111111101010","111111111111100100","000000000000000011","111111111111110110","000000000000001110","111111111111111111","111111111111100011","000000000000010010","111111111111110011","111111111111101001","111111111111101001","000000000000011001","000000000000001100","000000000000100111","000000000000011010","000000000000001010","000000000000001010","111111111111111101","111111111111111011","111111111111110101","111111111111100100","111111111111110010","111111111111111111","111111111111110010","000000000000000110","000000000000010110","111111111111111000","000000000000001010","000000000000001010","111111111111101011","111111111111100100","000000000000000101","111111111111110010","111111111111101010","000000000000000000","000000000000001100","000000000000010100","111111111111111011","111111111111100101","111111111111101110","000000000000001001","000000000000011000","111111111111011111","000000000000011001","000000000000010111","111111111111111100","111111111111110011","000000000000000110","111111111111110100","111111111111111101","111111111111101110","000000000000000001","000000000000010011","111111111111010001","111111111111100010","111111111111101011","111111111111111010","111111111111101011","000000000000000101","111111111111110010","111111111111111111","000000000000001011","111111111111110011","111111111111101110","111111111111111111","111111111111101110","111111111111101100","000000000000000001","000000000000001010","000000000000000010","111111111111111010","111111111111110101","111111111111111010","111111111111101111","111111111111101111","111111111111110110","111111111111110101","111111111111110111","111111111111110001","111111111111111000","000000000000101111","000000000000010001","111111111111110110","111111111111111010","111111111111011011","000000000000011000","000000000000010100","000000000000000101"),
("000000000000000110","000000000000100111","000000000000001110","000000000000000000","000000000000101000","111111111111110000","111111111111011010","111111111111110111","111111111111101001","000000000000000111","000000000000001000","000000000000000101","111111111111111101","000000000000100111","111111111111100010","111111111111101010","000000000000001011","111111111111101000","000000000000000001","000000000000000000","000000000000001110","111111111111101111","111111111111100101","111111111111111001","111111111111110011","111111111111111110","000000000000010011","111111111111111000","000000000000000100","000000000000001011","000000000000000100","000000000000011000","111111111111101101","000000000000000011","000000000000001100","000000000000000111","000000000000000011","000000000000001110","000000000000010100","000000000000010001","111111111111111111","000000000000100000","111111111111011111","000000000000001101","111111111111110101","000000000000010000","111111111111100011","000000000000110100","111111111111111000","111111111111010111","111111111111101011","111111111111111010","111111111111111101","111111111111111101","000000000000010000","111111111111100010","111111111111111110","111111111111100000","111111111111100100","000000000000001011","111111111111111001","111111111111111010","111111111111100001","111111111111111000","000000000000010110","000000000000000100","111111111111100110","111111111111101100","000000000000010011","111111111111111011","111111111111101001","000000000000000011","000000000000011000","111111111111101110","111111111111111000","000000000000010010","000000000000000001","111111111111011001","111111111111100000","111111111111100011","000000000000000010","111111111111111000","000000000000000000","000000000000011010","000000000000011110","000000000000010010","000000000000001001","000000000000100100","111111111111110011","000000000000001101","000000000000010000","111111111111011010","000000000000000001","111111111111111011","111111111111010110","111111111111101010","000000000000010000","111111111111100000","000000000000101110","111111111111110100","111111111111100001","000000000000001101","111111111111011111","111111111111100011","000000000000000111","111111111111010001","111111111111100110","111111111111010100","000000000000011000","111111111111101111","111111111111100111","111111111111101010","111111111111011101","111111111111110010","111111111111101111","000000000000000001","111111111111011010","000000000000100011","000000000000001100","000000000000011100","000000000000100110","000000000000100011","000000000000000010","000000000000000101","000000000000010001","000000000000001001","111111111111011011","000000000000010110"),
("111111111111101110","000000000000000000","111111111111101100","000000000000001000","111111111111101100","000000000000010000","000000000000000000","000000000000000110","111111111111110000","111111111111111100","111111111111110110","000000000000001001","000000000000001010","111111111111110110","000000000000000001","111111111111110111","000000000000010010","000000000000000011","000000000000000000","000000000000000101","000000000000010010","111111111111101100","000000000000000000","111111111111111110","000000000000001111","111111111111111010","000000000000010000","000000000000000011","000000000000010100","111111111111110011","111111111111111000","000000000000010010","000000000000000011","111111111111110101","111111111111101110","000000000000001101","111111111111111000","000000000000010001","111111111111111111","111111111111111000","111111111111110010","111111111111110010","000000000000000000","000000000000000000","111111111111111000","000000000000001111","000000000000010011","111111111111111110","000000000000000011","000000000000010000","000000000000000001","000000000000010011","111111111111101100","000000000000001001","000000000000001110","111111111111110010","000000000000001111","111111111111110110","000000000000000000","111111111111111100","000000000000010000","000000000000000111","111111111111111011","111111111111110000","111111111111111110","111111111111111110","000000000000000101","111111111111110011","000000000000000000","111111111111101101","111111111111101101","111111111111110100","000000000000001011","000000000000010010","111111111111111001","111111111111111011","111111111111110110","111111111111111101","000000000000000000","000000000000001110","000000000000001010","111111111111111110","000000000000001111","000000000000010001","000000000000001010","111111111111110000","000000000000000101","111111111111111110","111111111111101111","000000000000001011","000000000000000100","111111111111110001","000000000000000000","111111111111110110","111111111111111011","111111111111110011","111111111111110001","111111111111111100","111111111111101101","000000000000000001","000000000000010001","000000000000001010","000000000000010000","111111111111101101","000000000000000101","000000000000001110","000000000000001100","000000000000000101","000000000000001001","000000000000000111","000000000000000001","111111111111110011","000000000000000110","111111111111110010","111111111111101110","111111111111110011","111111111111110111","000000000000000100","111111111111111011","000000000000001110","000000000000010001","000000000000001010","000000000000000011","111111111111111110","111111111111111110","000000000000000000","000000000000000111","000000000000010011"),
("111111111111111010","111111111111111000","000000000000001000","111111111111111010","000000000000010010","111111111111111011","000000000000001001","000000000000001101","000000000000010000","000000000000001110","000000000000000011","000000000000000100","000000000000000000","111111111111111110","000000000000000111","111111111111110110","000000000000001001","000000000000010011","000000000000000011","111111111111101100","111111111111111010","111111111111110010","111111111111111100","000000000000001110","111111111111110100","000000000000000110","111111111111111010","000000000000000101","000000000000000100","111111111111110101","111111111111110110","111111111111110111","000000000000010001","000000000000010011","111111111111111110","111111111111111101","000000000000001111","111111111111101111","000000000000001110","111111111111101110","000000000000010011","000000000000000111","000000000000010011","111111111111110000","000000000000001011","000000000000000000","111111111111111100","111111111111111000","000000000000000000","000000000000000011","000000000000000100","000000000000000010","111111111111110101","000000000000000000","111111111111101111","111111111111110001","111111111111111110","000000000000010000","000000000000000000","000000000000010010","000000000000000011","000000000000000101","111111111111111010","000000000000010000","000000000000001001","111111111111111010","000000000000010001","000000000000000010","000000000000000010","000000000000010100","111111111111111011","111111111111111010","000000000000000001","111111111111110111","000000000000000110","000000000000000100","000000000000001110","111111111111101110","000000000000010011","000000000000001111","111111111111110010","111111111111101101","111111111111111000","111111111111111000","000000000000010100","111111111111110101","000000000000000010","111111111111110001","000000000000010010","000000000000000010","000000000000010010","111111111111111111","111111111111110101","000000000000000100","111111111111110111","000000000000001100","111111111111110110","000000000000001110","111111111111111101","000000000000000110","000000000000010000","111111111111101100","000000000000001101","000000000000001111","000000000000000111","111111111111111001","111111111111110000","111111111111110000","111111111111110100","111111111111101100","111111111111111100","111111111111111111","111111111111111010","000000000000000101","000000000000000101","000000000000000111","111111111111101101","000000000000000011","000000000000010100","000000000000000001","111111111111110110","000000000000010000","000000000000001010","111111111111101100","000000000000000011","000000000000000011","000000000000001001","000000000000001100"),
("000000000000000010","111111111111111101","000000000000010010","111111111111111011","111111111111101110","000000000000010000","000000000000000000","000000000000000011","000000000000001010","000000000000001011","111111111111101101","000000000000010100","111111111111111011","111111111111111111","000000000000010011","000000000000000110","111111111111110000","111111111111110001","111111111111101100","111111111111111011","111111111111110010","111111111111110011","111111111111110011","000000000000000001","111111111111111011","111111111111111011","111111111111110101","000000000000001101","111111111111111110","000000000000000011","111111111111111010","111111111111101110","000000000000000110","000000000000001000","000000000000000100","000000000000000100","111111111111110000","111111111111111111","000000000000000110","111111111111111111","000000000000000101","000000000000010010","000000000000000001","000000000000001101","111111111111110101","111111111111110111","000000000000001111","000000000000001011","111111111111110001","111111111111111001","000000000000000111","111111111111111110","111111111111111010","000000000000001011","000000000000010100","000000000000001010","000000000000001110","111111111111101101","000000000000001011","111111111111110110","111111111111111011","111111111111111101","000000000000001110","111111111111101110","111111111111110010","000000000000010100","000000000000001011","111111111111111000","111111111111111001","111111111111111011","111111111111111111","000000000000001010","000000000000000011","000000000000001011","111111111111110010","000000000000001000","000000000000001101","111111111111110000","111111111111111111","111111111111110101","111111111111101111","111111111111110010","000000000000001001","111111111111101110","000000000000000011","000000000000000101","111111111111110111","000000000000001001","111111111111110010","111111111111101101","000000000000000000","000000000000001101","000000000000010010","111111111111111110","111111111111111100","111111111111111111","000000000000000101","000000000000001111","000000000000000010","000000000000000001","111111111111111101","111111111111111110","111111111111101100","000000000000001011","000000000000001110","111111111111110010","000000000000000000","000000000000000000","111111111111110101","000000000000010000","000000000000001110","111111111111110100","000000000000001101","111111111111110001","111111111111101100","111111111111110100","111111111111111111","000000000000000100","111111111111101101","111111111111110000","111111111111101111","000000000000000101","111111111111101101","111111111111111111","111111111111101110","000000000000000001","111111111111111110","000000000000000011"),
("111111111111110001","000000000000000111","111111111111111111","111111111111101110","000000000000001111","000000000000000000","111111111111101000","000000000000011110","000000000000000111","000000000000001101","000000000000001100","000000000000000010","111111111111110010","000000000000000000","111111111111110110","111111111111101100","111111111111111111","111111111111110110","000000000000010110","111111111111111100","111111111111100111","111111111111111100","000000000000000101","111111111111010110","000000000000000100","000000000000001011","000000000000000001","000000000000000111","000000000000101010","000000000000010110","111111111111100000","000000000000101001","000000000000010011","000000000000000010","000000000000000010","000000000000100100","111111111111111000","000000000000010111","000000000000100100","000000000000110110","000000000000011110","111111111111100101","111111111111111000","111111111111100000","111111111111111001","000000000000010001","111111111111111101","111111111111110101","000000000000010111","000000000000100000","000000000000100000","000000000000010011","111111111111110101","000000000000100010","000000000000010011","000000000000001001","000000000000001110","000000000000000011","111111111111110001","111111111111111110","000000000000001011","000000000000000001","000000000000001000","000000000000001110","111111111111101110","111111111111110000","111111111111011000","111111111111110111","000000000000001101","111111111111110100","000000000000010001","000000000000101001","000000000000011101","000000000000000010","111111111111111111","111111111111110111","111111111111110101","111111111111110111","111111111111100111","111111111111111101","111111111111110010","000000000000000111","000000000000010100","000000000000011110","111111111111111000","000000000000000000","111111111111101100","000000000000010111","111111111111111100","000000000000000100","111111111111101010","000000000000011011","000000000000100010","111111111111110110","111111111111100101","000000000000010110","111111111111110000","111111111111101000","000000000000000101","000000000000001001","111111111111101010","111111111111101010","000000000000001000","000000000000001000","000000000000000100","111111111111110100","111111111111101011","000000000000001000","000000000000010101","000000000000000100","000000000000000000","111111111111101110","000000000000001000","000000000000010001","000000000000110101","111111111111111001","000000000000001010","000000000000000011","000000000000000001","111111111111111100","111111111111110010","111111111111010010","111111111111110100","000000000000001000","111111111111100110","111111111111111111","111111111111111101","000000000000010101"),
("111111111111111001","000000000000001111","111111111111111110","111111111111010101","111111111111100001","111111111111001110","111111111111100100","000000000000011010","111111111111100000","111111111111111000","111111111111010111","000000000000110100","111111111111000101","111111111111111110","000000000000000011","111111111111110101","000000000000110100","111111111111010010","000000000000010001","000000000000010001","111111111111100001","111111111111110011","111111111111110110","111111111111100111","111111111111110001","111111111111100101","111111111111110100","111111111111111001","000000000000000000","000000000000010101","111111111111110001","000000000000011001","000000000000101100","000000000000010111","111111111111011001","111111111111110101","000000000000000010","000000000000010010","000000000000100111","000000000000111111","000000000000011010","111111111111010110","111111111111100111","111111111111100001","000000000000011101","000000000000000101","111111111111101110","111111111111100001","000000000000111010","000000000000001110","111111111111111101","111111111111111011","111111111111111100","000000000000100111","000000000000100010","111111111111010010","000000000000100101","000000000000010011","000000000000000000","111111111111110111","000000000000010110","000000000000011101","111111111111101111","111111111111101111","111111111111111000","000000000000000111","111111111111011101","000000000000000000","000000000000101011","000000000000000011","000000000000001001","000000000000101011","000000000000011000","111111111111110111","000000000000100011","111111111111111010","111111111111111101","000000000000001110","111111111111011000","000000000000011000","111111111111111101","111111111111111110","111111111111110101","000000000000101110","000000000000001000","000000000000001000","000000000000001011","000000000000101110","000000000000001001","000000000000010000","111111111111101000","000000000000000001","000000000000001101","111111111111100011","111111111111110001","000000000000001101","000000000000000000","000000000000000101","000000000000100011","000000000000000101","111111111111110010","000000000000011011","000000000000000011","000000000000000010","111111111111010111","111111111111110111","111111111111111100","000000000000001110","000000000000100101","111111111111100000","000000000000000000","111111111111110001","000000000000001101","000000000000100101","000000000000001010","000000000000000001","000000000000100000","000000000000101101","111111111111100001","000000000000010101","111111111111111101","111111111111100010","111111111111101011","111111111111101110","111111111111100011","000000000000001000","111111111111111000","000000000000010101"),
("111111111111011100","111111111111100110","000000000000000011","111111111111010101","111111111111110000","111111111111011000","111111111111111000","111111111111111011","000000000000001101","000000000000010100","111111111111000101","000000000000011001","000000000000001110","000000000000001100","111111111111111011","111111111111100110","000000000000000001","111111111111010101","111111111111110000","000000000000111001","000000000000000001","000000000000000000","000000000000011000","111111111111010100","111111111111100010","111111111111100100","111111111111100000","111111111111111111","000000000000011000","000000000000000110","111111111111100011","000000000000011110","000000000000010011","000000000000000110","111111111111110100","111111111111111010","000000000000010011","000000000000001110","000000000000011000","000000000000111101","000000000000100100","111111111111110111","000000000000001011","111111111111001111","111111111111111111","000000000000000001","111111111111010000","000000000000001000","000000000000011011","000000000000110001","000000000000001111","000000000000000010","111111111111101011","000000000000000110","000000000000100000","111111111111101111","000000000000001101","000000000000011010","000000000000010101","000000000000000000","000000000000010001","000000000000100111","111111111111110001","111111111111010001","111111111111101001","000000000000001000","111111111111001111","000000000000100000","000000000000111011","111111111111011101","111111111111111100","000000000000000110","000000000000100110","000000000000010101","000000000000011100","000000000000110100","111111111111101001","000000000000001010","111111111111101111","111111111111111010","111111111111111110","111111111111111000","000000000000000001","000000000000101001","111111111111101111","000000000000011111","111111111111111111","000000000000100011","000000000000100100","000000000000101011","000000000000001101","000000000000001110","000000000000010111","111111111111101010","111111111111111110","000000000000011110","000000000000001111","000000000000001101","000000000000000010","000000000000100011","111111111111101110","111111111111101100","000000000000010111","111111111111100100","111111111111100010","111111111111101011","111111111111110011","111111111111111001","000000000000011110","111111111111101010","111111111111111011","111111111111010101","000000000000001101","000000000000100001","000000000000010100","111111111111111101","000000000000010111","000000000000111101","000000000000000011","000000000000101000","000000000000011110","111111111111111010","111111111111110110","111111111111111100","111111111111101111","111111111111110111","111111111111111111","000000000000011011"),
("111111111111111101","111111111111100001","000000000000001110","111111111111100000","111111111111101100","111111111111010111","111111111111110111","000000000000000111","111111111111101101","000000000000001101","111111111111011101","000000000000001110","000000000000000010","000000000000001011","111111111111110001","111111111111111101","111111111111010100","111111111111101111","111111111111101110","000000000000000100","000000000000010000","000000000001000011","111111111111111001","000000000000000000","000000000000000000","111111111111010101","111111111111011111","000000000000001100","000000000000000101","000000000000000010","111111111111101001","000000000000010100","111111111111111001","111111111111111110","111111111111111011","111111111111110100","000000000000100001","111111111111110101","000000000000010111","000000000000001001","000000000000001111","000000000000000100","111111111111110110","111111111111011101","111111111111111101","000000000000001110","111111111111110000","000000000000010111","000000000000001111","000000000000011110","000000000000000000","111111111111101110","000000000000000010","000000000000010011","000000000000011111","111111111111110001","000000000000000011","000000000000101111","000000000000100010","000000000000001110","000000000000101100","000000000000000010","111111111111101011","111111111111001111","111111111111011110","000000000000010010","000000000000000100","000000000000000111","000000000000010100","111111111111111011","111111111111100101","000000000000000101","000000000000000100","000000000000010000","000000000000001011","000000000000100101","111111111111011001","000000000000010111","000000000000001001","111111111111110100","111111111111101100","111111111111110001","111111111111101110","000000000000011000","111111111111100010","000000000000010101","000000000000011010","000000000000000110","111111111111110100","000000000000000000","000000000000000111","000000000000000111","111111111111100001","111111111111110100","000000000000011100","000000000000100011","000000000000000100","000000000000010100","111111111111100011","000000000000100100","111111111111100011","111111111111111001","000000000000011011","111111111111010011","111111111111011111","111111111111011001","000000000000000001","000000000000011011","000000000000010000","111111111111110110","000000000000001110","111111111111111101","111111111111110110","000000000000001110","111111111111110000","111111111111110101","000000000000001110","000000000000011001","111111111111111000","000000000000101101","000000000000010111","000000000000000110","111111111111101101","111111111111100111","000000000000000000","111111111111101000","000000000000000111","000000000000001101"),
("111111111111111001","111111111111101101","111111111111110100","111111111111110100","111111111111001010","111111111111011010","111111111111110000","111111111111010110","000000000000000111","111111111111111101","111111111111101011","000000000000010111","111111111111110111","000000000000000100","111111111111000000","111111111111110100","111111111111110011","111111111111111010","000000000000000000","000000000000001100","111111111111111110","000000000000111001","111111111111110010","111111111111110011","111111111111101101","111111111111100001","111111111111001111","111111111111011001","000000000000011110","000000000000000010","111111111111011111","000000000000000011","000000000000001000","111111111111100100","111111111111101010","111111111111111110","000000000000000000","111111111111111111","000000000000100101","000000000000001001","000000000000001011","000000000000010000","111111111111111010","111111111111000100","111111111111110010","000000000000011101","111111111111011111","111111111111101111","000000000000001011","000000000000101000","000000000000001111","111111111111101011","000000000000000001","111111111111110010","000000000000101001","000000000000010100","111111111111101011","000000000000011011","000000000000010101","000000000000001100","111111111111111010","000000000000000010","111111111111111101","111111111111101100","111111111110111000","000000000000010111","111111111111010010","111111111111111101","000000000000011110","000000000000001110","111111111111100011","111111111111111101","111111111111011010","000000000000001110","000000000000010111","000000000000011010","111111111111100011","000000000000000010","000000000000000011","000000000000011000","111111111111101110","111111111111111010","111111111111111010","000000000000100101","111111111111110111","000000000000001001","000000000000011000","000000000000100000","000000000000001101","000000000000000000","000000000000010101","000000000000010111","111111111111000110","111111111111110110","111111111111110100","000000000000000100","111111111111110101","000000000000000000","111111111111011101","000000000000100011","111111111111101000","000000000000000101","111111111111111100","111111111111111001","111111111111110000","111111111111101011","000000000000001101","000000000000001000","000000000000100111","111111111111110101","000000000000010011","111111111111111100","111111111111111101","000000000000000101","000000000000011010","000000000000000010","111111111111111000","000000000000010111","000000000000000000","000000000000011011","000000000000001010","111111111111110000","111111111111101001","000000000000011111","000000000000000010","111111111111101100","111111111111110011","000000000000001010"),
("111111111111111000","111111111111100110","111111111111110011","111111111111011101","111111111111101000","111111111111101101","000000000000000001","111111111111111111","000000000000010011","111111111111111110","111111111111010111","000000000000000001","000000000000001001","000000000000000111","111111111111010101","111111111111101001","000000000000000000","111111111111100101","111111111111111010","000000000000100101","000000000000000100","000000000000101001","111111111111101011","000000000000001000","000000000000000011","111111111111101101","111111111111010101","111111111111110001","000000000000100010","000000000000001000","111111111111101001","000000000000000011","000000000000000101","111111111111100011","111111111111111111","111111111111101110","000000000000000000","111111111111100110","000000000000010010","000000000000000000","000000000000000011","000000000000001010","111111111111011100","111111111111001000","000000000000010101","000000000000000000","111111111110111110","111111111111010011","000000000000010010","000000000000011101","000000000000000000","000000000000001000","000000000000011100","000000000000000100","000000000000010010","000000000000100100","000000000000001011","000000000000100001","000000000000100100","000000000000010000","111111111111111001","111111111111111010","111111111111111101","111111111111011110","111111111111101001","000000000000001010","111111111111110111","111111111111101001","000000000000110111","000000000000000101","000000000000000000","111111111111110110","111111111110111100","111111111111111010","000000000000001001","000000000000100111","111111111111111100","000000000000010001","000000000000011110","000000000000000101","111111111111100111","000000000000010001","111111111111110111","000000000000000110","000000000000000000","000000000000011000","000000000000011001","000000000000100011","000000000000000001","111111111111110100","000000000000001000","000000000000010111","111111111111100000","111111111111101110","111111111111101010","000000000000011111","000000000000000000","000000000000000100","111111111111110000","000000000000010001","111111111111011110","111111111111100100","000000000000001011","111111111111101100","111111111111101100","111111111111101110","000000000000000100","111111111111111111","000000000000011101","111111111111110100","000000000000010101","000000000000000000","111111111111110000","000000000000001001","000000000000000000","000000000000001101","000000000000010010","111111111111111101","000000000000011000","000000000000001101","000000000000011000","000000000000001011","111111111111100010","111111111111111100","000000000000000110","111111111111110100","000000000000001000","000000000000010110"),
("000000000000010000","111111111111011101","000000000000000000","111111111111110111","111111111111110001","111111111111111101","000000000000000010","111111111111101101","000000000000000000","000000000000000100","111111111111101101","000000000000010101","111111111111110011","000000000000100111","111111111111010101","000000000000000011","000000000000000001","111111111111110110","111111111111110110","000000000000010011","000000000000001011","000000000001001001","000000000000001011","000000000000000001","000000000000000000","111111111111110011","111111111111101111","111111111111100101","000000000000000110","111111111111101101","111111111111101100","111111111111111000","000000000000001000","111111111111111100","111111111111101101","000000000000000001","000000000000010011","111111111111110111","000000000000000101","111111111111101010","000000000000000000","000000000000010111","111111111110111101","111111111110111001","000000000000011111","000000000000000111","111111111111001010","111111111111111010","000000000000000111","000000000000001001","111111111111111110","000000000000010011","000000000000001101","111111111111111111","111111111111111011","000000000000000011","111111111111110100","000000000000000111","000000000000000001","111111111111101101","000000000000010010","000000000000010010","111111111111110000","000000000000010000","000000000000000010","000000000000000000","111111111111111001","000000000000001010","000000000000011001","111111111111111011","000000000000001101","000000000000010011","111111111111000111","111111111111110101","111111111111100100","000000000000101100","000000000000000110","111111111111111111","111111111111110011","111111111111111110","000000000000000001","111111111111110101","000000000000000000","111111111111101100","000000000000010001","111111111111101101","000000000000010110","111111111111111001","000000000000000111","000000000000010111","000000000000001111","000000000000100101","111111111111101000","111111111111110000","111111111111100100","000000000000100001","000000000000001101","000000000000001011","111111111111111110","111111111111111100","111111111111101010","111111111111100010","000000000000010100","000000000000100100","111111111111111110","111111111111111111","000000000000000100","111111111111110110","000000000000001101","111111111111110110","000000000000011001","000000000000010000","000000000000010010","000000000000001110","111111111111111011","000000000000001101","000000000000001111","000000000000011001","000000000000010101","000000000000001100","000000000000100101","000000000000000100","111111111111110101","000000000000011010","111111111111100010","111111111111111111","000000000000010001","000000000000000010"),
("111111111111111000","111111111111101001","111111111111111100","000000000000001001","000000000000000001","111111111111101110","000000000000000100","000000000000000100","111111111111101101","000000000000000101","000000000000000000","000000000000110001","111111111111011101","000000000000010011","111111111111111011","000000000000010100","111111111111011011","000000000000001110","000000000000000010","000000000000010010","111111111111101001","000000000000011111","111111111111110011","111111111111111110","000000000000001111","111111111111110100","111111111111111101","111111111111110101","000000000000010100","000000000000001111","111111111111100100","111111111111101010","000000000000001000","111111111111111111","000000000000001100","111111111111111100","111111111111101110","000000000000010000","000000000000101011","111111111111110000","000000000000000100","000000000000011011","111111111110101000","111111111111011000","111111111111111111","000000000000010111","111111111111100011","000000000000000000","000000000000100010","111111111111101110","000000000000000111","000000000000001111","000000000000001100","111111111111100001","000000000000010000","000000000000010010","111111111111110111","000000000000001110","111111111111110001","000000000000001001","000000000000000011","000000000000000110","000000000000010010","000000000000001000","111111111111101011","000000000000001111","000000000000000101","111111111111111110","000000000000011110","000000000000000011","000000000000000000","000000000000010011","111111111111010111","111111111111100010","000000000000000000","000000000000101111","000000000000000011","000000000000001011","000000000000000110","000000000000000000","000000000000000010","000000000000000011","111111111111001100","111111111111110001","000000000000011010","111111111111101110","000000000000011110","000000000000011101","000000000000000100","000000000000000111","111111111111110100","000000000000001110","111111111111111001","111111111111111110","111111111111101101","000000000000001011","000000000000111010","000000000000000110","111111111111111110","000000000000000010","111111111111111010","111111111111111001","000000000000010011","000000000000001101","000000000000001000","111111111111110110","000000000000010110","111111111111101001","111111111111110110","111111111111110100","000000000000000011","111111111111111110","000000000000000110","000000000000011100","111111111111110111","000000000000001101","111111111111100101","000000000000100001","000000000000011101","111111111111111100","000000000000010001","000000000000100110","111111111111010111","111111111111110010","000000000000001110","111111111111110101","000000000000000011","111111111111111001"),
("111111111111100011","111111111111110000","000000000000000001","111111111111111111","111111111111001011","111111111111100100","000000000000001111","111111111111111001","000000000000010011","111111111111110010","000000000000001110","000000000000010111","111111111111011110","111111111111111000","111111111111111110","111111111111111110","111111111111110101","000000000000000010","000000000000000000","111111111111111110","000000000000000000","000000000000001010","000000000000000111","000000000000001001","111111111111111110","000000000000000111","000000000000010001","000000000000000000","111111111111111010","000000000000001000","000000000000001011","111111111111111011","000000000000010101","111111111111110101","000000000000001110","111111111111111010","111111111111100111","000000000000010010","000000000000010110","111111111111111101","000000000000011110","111111111111111000","111111111111001110","000000000000000001","000000000000011001","000000000000000010","111111111111011011","111111111111101111","000000000000010010","000000000000001010","000000000000010110","000000000000010000","000000000000011010","111111111111110001","111111111111110100","111111111111111010","000000000000010110","111111111111111110","111111111111111011","000000000000010000","000000000000001001","111111111111111001","111111111111111101","111111111111111000","111111111111110011","111111111111110110","000000000000000001","000000000000000000","000000000000010110","000000000000000011","000000000000001001","111111111111110111","111111111111110011","000000000000001000","111111111111111001","000000000000011010","000000000000000010","000000000000001110","000000000000001010","111111111111110001","000000000000001010","000000000000000000","111111111111001010","111111111111101111","000000000000000110","000000000000001000","000000000000000100","000000000000000101","111111111111101010","000000000000000111","000000000000001010","000000000000100000","000000000000001000","000000000000001100","111111111111100011","000000000000001011","000000000000101101","111111111111111100","111111111111110000","000000000000011001","111111111111111101","111111111111110101","000000000000010100","000000000000000111","000000000000000110","000000000000000101","000000000000100001","000000000000000001","000000000000010011","111111111111110000","000000000000001001","000000000000001101","000000000000001001","111111111111111101","111111111111110111","111111111111110101","111111111111111011","111111111111111111","000000000000001001","111111111111111011","000000000000000010","000000000000000010","111111111111100101","111111111111011010","111111111111110101","111111111111101011","000000000000000010","000000000000011100"),
("111111111111011110","111111111111010010","000000000000100101","111111111111110101","111111111111101110","111111111111011111","000000000000011101","111111111111110101","111111111111110010","000000000000000110","111111111111111100","000000000000100101","000000000000000100","111111111111100100","111111111111111111","111111111111111011","111111111111111100","000000000000010101","111111111111110101","000000000000000101","000000000000000010","111111111111100000","111111111111111101","000000000000000110","000000000000001110","000000000000001010","000000000000100000","111111111111111111","000000000000001100","000000000000010000","000000000000000100","000000000000000110","111111111111111111","111111111111110111","000000000000000100","000000000000000001","000000000000000000","000000000000011100","000000000000000010","111111111111111011","111111111111111010","000000000000000101","111111111111010001","111111111111101100","000000000000001111","000000000000001011","111111111111110010","111111111111110100","000000000000100000","111111111111111010","111111111111111001","000000000000001001","000000000000010111","111111111111111001","111111111111111110","000000000000101001","000000000000000010","000000000000000111","000000000000010101","111111111111110011","000000000000001110","111111111111110100","000000000000100010","000000000000000110","111111111111100101","000000000000001101","000000000000001011","000000000000000000","000000000000010010","000000000000001100","000000000000000101","000000000000011000","111111111111011001","111111111111110010","111111111111101011","000000000000010100","000000000000000011","111111111111111110","111111111111111000","111111111111110101","000000000000000010","000000000000010101","111111111111011111","000000000000010010","000000000000011000","111111111111111001","000000000000001001","111111111111111010","111111111111110000","000000000000001101","111111111111101011","000000000000010101","000000000000000000","111111111111101010","111111111111111001","000000000000010000","000000000000010100","000000000000001011","000000000000000001","000000000000100000","111111111111100010","111111111111111011","000000000000001101","000000000000100011","000000000000000001","000000000000001000","000000000000100010","000000000000011011","000000000000000110","111111111111100111","000000000000100001","000000000000100001","000000000000000110","000000000000000011","000000000000011000","111111111111101000","111111111111111001","111111111111111011","000000000000010001","111111111111111110","000000000000001101","000000000000000110","000000000000000111","111111111111110101","111111111111110110","111111111111111010","000000000000001110","000000000000000111"),
("111111111111110010","111111111111111000","000000000000000000","000000000000011101","111111111111101011","111111111111011101","000000000000001100","111111111111110100","000000000000000110","000000000000001101","000000000000010011","000000000000101000","000000000000000000","111111111111011100","000000000000000101","000000000000001001","000000000000000001","000000000000010001","000000000000001000","000000000000001000","000000000000010111","111111111111010110","000000000000000111","000000000000010100","000000000000001111","000000000000010100","000000000000010000","111111111111110110","000000000000001001","000000000000011011","000000000000001000","111111111111111010","000000000000100110","111111111111101111","111111111111110111","111111111111110010","000000000000001101","000000000000000011","111111111111110111","000000000000000111","000000000000011001","111111111111111011","111111111111101010","000000000000001100","000000000000011011","000000000000000101","111111111111110001","111111111111100111","000000000000010100","111111111111111101","000000000000001011","000000000000001110","000000000000000111","111111111111101010","111111111111011011","111111111111110010","000000000000100010","000000000000010010","000000000000010110","111111111111111111","000000000000100011","111111111111111110","000000000000100111","000000000000000111","111111111111101101","000000000000001101","000000000000001111","111111111111100110","000000000000000000","111111111111111010","111111111111111111","000000000000011011","111111111111110001","111111111111111011","111111111111110101","111111111111101100","000000000000000011","111111111111111010","111111111111101011","000000000000001100","111111111111101100","000000000000000101","111111111111011000","000000000000001110","000000000000011010","111111111111101101","000000000000100100","000000000000000100","000000000000000010","000000000000000000","111111111111010101","000000000000001100","111111111111110101","111111111111101101","111111111111111011","000000000000000000","000000000000010111","000000000000001100","111111111111110100","111111111111111011","111111111111100111","000000000000010000","000000000000001000","000000000000001001","000000000000101010","000000000000010001","111111111111111111","000000000000011111","111111111111100010","000000000000000001","000000000000001101","000000000000011101","000000000000100000","000000000000001010","111111111111111110","000000000000001110","000000000000010101","000000000000000011","000000000000011010","111111111111111010","000000000000001010","000000000000001010","111111111111110101","111111111111110110","111111111111101010","000000000000011011","000000000000011100","000000000000001001"),
("000000000000001001","000000000000000000","000000000000000111","000000000000011101","111111111111101010","111111111111011011","000000000000010000","000000000000001001","111111111111111000","000000000000011011","000000000000010100","000000000001001000","111111111111100010","111111111111010010","000000000000000100","000000000000011011","111111111111101000","000000000000010000","000000000000011101","000000000000010001","000000000000000011","111111111111101101","111111111111100100","000000000000101000","000000000000101000","111111111111101110","000000000000101110","111111111111110100","000000000000001010","000000000000011001","000000000000001000","111111111111011101","000000000000011011","111111111111111000","000000000000000110","000000000000000110","111111111111111011","000000000000010111","111111111111111100","000000000000010000","111111111111111111","111111111111110100","111111111111111100","111111111111110001","000000000000010111","000000000000001100","111111111111110101","111111111111110011","000000000000100010","000000000000010110","000000000000000000","000000000000010101","000000000000000110","111111111111111111","111111111111111111","111111111111110110","000000000000010001","000000000000000010","000000000000000101","111111111111111000","000000000000000111","111111111111110100","000000000000010100","111111111111101011","111111111111111010","000000000000010100","111111111111110110","111111111111101111","000000000000000111","000000000000011010","111111111111111110","000000000000011101","000000000000000000","111111111111111010","111111111111100010","111111111111110101","111111111111110100","000000000000010001","111111111111101100","000000000000000001","000000000000000010","000000000000001110","111111111111011011","111111111111111101","000000000000001111","000000000000000000","000000000000011101","000000000000001100","000000000000000111","111111111111101010","111111111111110001","000000000000011100","111111111111111111","111111111111101111","111111111111111100","000000000000010010","000000000000010011","000000000000001110","111111111111100100","111111111111110001","111111111111100000","000000000000000010","000000000000001111","000000000000000101","000000000000011111","000000000000001110","000000000000000100","000000000000000111","111111111111101011","111111111111111100","111111111111110110","000000000000010011","000000000000100001","000000000000010011","000000000000011111","111111111111101100","000000000000000100","111111111111110101","111111111111111110","000000000000010110","000000000000011101","000000000000011100","000000000000000001","111111111111110001","111111111111110110","000000000000000100","000000000000001010","000000000000001000"),
("000000000000001101","000000000000100000","111111111111111110","000000000000001111","111111111111111011","111111111111010101","000000000000000011","000000000000100000","111111111111111100","000000000000010000","000000000000100010","000000000000110110","111111111111111000","000000000000000000","111111111111110010","000000000000101100","111111111111100100","000000000000001110","000000000000100011","000000000000001111","111111111111100101","111111111111110111","111111111111110001","000000000000001011","000000000000011111","111111111111111010","000000000000011011","000000000000001011","000000000000001110","000000000000010111","000000000000000100","111111111111110001","000000000000100010","000000000000000000","000000000000010101","000000000000001110","111111111111111001","000000000000000110","111111111111110010","000000000000011011","111111111111111101","000000000000010001","111111111111111110","111111111111110010","000000000000100001","111111111111111101","000000000000000111","111111111111111101","000000000000001111","000000000000010010","000000000000010001","000000000000010011","111111111111111011","111111111111100001","111111111111111011","000000000000000101","111111111111111101","000000000000000000","000000000000000110","000000000000000000","000000000000000011","000000000000011000","000000000000000111","000000000000000000","000000000000000000","111111111111111000","111111111111010111","111111111111101101","000000000000011001","000000000000001010","000000000000001101","000000000000010011","111111111111100100","000000000000010101","111111111111010101","111111111111111011","000000000000001011","000000000000000110","111111111111100110","111111111111111111","000000000000001100","000000000000000000","111111111111100000","111111111111110110","000000000000100001","111111111111111001","000000000000101111","000000000000001110","000000000000010001","000000000000000000","000000000000000100","000000000000010001","000000000000000111","111111111111101000","111111111111110111","000000000000001000","000000000000001010","000000000000011000","111111111111101111","111111111111101010","111111111111111010","000000000000000010","111111111111111000","000000000000000011","000000000000000000","000000000000010010","000000000000000000","000000000000100001","111111111111010010","111111111111111000","000000000000000000","000000000000000001","000000000000001100","000000000000100000","000000000000011010","111111111111101011","000000000000001110","000000000000011010","000000000000001000","000000000000010001","000000000000011110","111111111111101111","111111111111111011","000000000000001111","111111111111100111","000000000000010011","000000000000001001","111111111111111001"),
("111111111111111111","000000000000100000","000000000000010001","000000000000010111","111111111111110100","111111111111101100","111111111111111110","000000000000010110","111111111111110010","000000000000001011","000000000000000001","000000000000011010","000000000000001011","111111111111100101","111111111111111010","000000000000011100","111111111111010111","000000000000000000","000000000000010011","000000000000001011","111111111111110110","000000000000000011","000000000000011110","000000000000000011","000000000000010010","000000000000001110","000000000000010101","000000000000000110","000000000000000001","000000000000000111","000000000000001011","111111111111110010","000000000000001000","000000000000001011","111111111111111011","111111111111110111","111111111111110100","000000000000000000","000000000000011010","000000000000001101","000000000000010001","111111111111111111","111111111111111111","000000000000000110","000000000000010000","111111111111010111","000000000000001111","111111111111111110","000000000000011000","111111111111111101","000000000000001110","000000000000001010","111111111111111011","000000000000001000","111111111111100011","111111111111101001","000000000000011011","000000000000000110","111111111111111011","000000000000000011","111111111111110110","111111111111111001","111111111111110110","111111111111110110","000000000000000111","000000000000000100","111111111111010001","111111111111110111","000000000000000110","000000000000001011","111111111111111101","000000000000010011","111111111111111110","111111111111110100","111111111111101110","000000000000001100","000000000000000000","111111111111111010","111111111111101001","111111111111111000","000000000000010101","000000000000000101","111111111111010011","111111111111101100","000000000000001111","111111111111011011","000000000000010001","111111111111110011","000000000000010000","000000000000000100","000000000000001001","000000000000000010","000000000000001101","111111111111100111","000000000000010010","000000000000001110","111111111111111110","000000000000000010","111111111111001101","111111111111100111","111111111111101111","000000000000000001","111111111111101000","000000000000000010","000000000000010101","000000000000011010","111111111111110111","000000000000010100","111111111111100011","000000000000000111","000000000000010110","000000000000001101","000000000000100000","000000000000001110","000000000000001110","111111111111111000","000000000000100010","111111111111110100","111111111111111001","000000000000001001","000000000000011101","111111111111101101","000000000000000010","000000000000000100","111111111111110101","000000000000001011","000000000000100011","111111111111111000"),
("000000000000001111","000000000000011101","111111111111111111","000000000000010100","000000000000000011","000000000000000110","111111111111110000","000000000000011000","000000000000000011","111111111111111111","000000000000000101","000000000000101010","000000000000000001","111111111111101010","000000000000101000","000000000000010010","111111111111101011","111111111111111110","000000000000010101","000000000000000000","111111111111110001","000000000000010010","000000000000000001","111111111111111100","000000000000000000","000000000000011010","000000000000010101","000000000000010000","000000000000001010","111111111111101110","000000000000001001","111111111111111101","000000000000110010","111111111111100111","111111111111111101","000000000000001001","111111111111111000","111111111111101010","000000000000010110","000000000000010101","000000000000001111","111111111111101111","000000000000000011","111111111111110001","000000000000011011","111111111111010010","111111111111111101","111111111111110000","000000000000010001","000000000000010101","111111111111110111","000000000000001000","111111111111110110","111111111111110100","111111111111011110","000000000000001110","000000000000100011","000000000000010000","111111111111111010","000000000000010001","111111111111110000","000000000000000011","111111111111100101","111111111111111000","000000000000001010","000000000000100000","111111111111100001","111111111111110011","111111111111111110","111111111111111100","000000000000001011","111111111111111010","111111111111110010","000000000000001000","000000000000001111","111111111111111011","111111111111111110","000000000000001011","000000000000001001","000000000000010010","000000000000000011","000000000000011100","111111111111000100","111111111111100010","000000000000010111","111111111111111110","000000000000100000","111111111111101111","000000000000110011","111111111111111100","111111111111110111","000000000000000001","000000000000000110","111111111111011100","111111111111111010","111111111111101010","111111111111111100","000000000000101111","111111111111100101","111111111111001100","111111111111101000","000000000000011111","000000000000001000","000000000000100000","111111111111101010","000000000000000100","000000000000000000","000000000000110010","000000000000000000","000000000000011010","000000000000000101","111111111111111101","000000000000001011","000000000000010001","000000000000011010","111111111111110010","000000000000101111","111111111111111100","111111111111111000","000000000000001101","000000000000010000","111111111111110111","111111111111100001","000000000000011100","111111111111100010","000000000000001111","000000000000100000","111111111111110011"),
("111111111111110111","000000000000011110","000000000000000111","000000000000001001","000000000000011101","111111111111101111","111111111111101100","000000000000101111","000000000000000000","000000000000100101","000000000000100000","000000000000011110","000000000000001111","111111111111101011","000000000000001101","000000000000010111","111111111111101110","111111111111111110","111111111111111001","000000000000000001","000000000000000111","000000000000011101","000000000000010101","111111111111000011","111111111111110111","000000000000001001","111111111111111011","000000000000000000","000000000000000101","000000000000000110","000000000000010011","111111111111111000","000000000000101011","111111111111111001","111111111111111101","111111111111110111","000000000000000000","111111111111100100","111111111111111111","000000000000011111","000000000000010000","111111111111010000","000000000000001101","000000000000000011","000000000000001010","111111111111110111","111111111111111011","111111111111011101","000000000000000111","000000000000001001","111111111111100010","000000000000010001","111111111111100000","000000000000010100","111111111111110001","111111111111111101","000000000000000000","000000000000000111","111111111111100100","111111111111110110","111111111111110001","000000000000010110","111111111111011001","000000000000000000","111111111111111110","111111111111110111","111111111111011111","111111111111101011","000000000000010001","000000000000010001","000000000000000001","000000000000010001","000000000000001110","000000000000000011","000000000000000010","111111111111111010","000000000000010010","000000000000000101","111111111111101010","111111111111110000","000000000000001101","000000000000100100","111111111110110010","111111111111101000","000000000000001100","000000000000000000","000000000000001100","111111111111111011","111111111111111101","000000000000000111","000000000000010110","000000000000010010","000000000000001000","111111111111111101","111111111111111110","111111111111100101","111111111111110101","000000000000011110","111111111111100101","111111111111000010","111111111111011001","000000000000001001","111111111111101101","111111111111110110","111111111111011101","000000000000001111","111111111111110000","000000000000001011","111111111111101101","000000000000010100","111111111111101101","000000000000000110","111111111111111101","111111111111101010","111111111111111110","000000000000000100","000000000000000100","000000000000001111","111111111111110101","000000000000010101","000000000000001011","111111111111110110","111111111111110111","000000000000000111","111111111111101110","000000000000001100","000000000000010011","000000000000010000"),
("000000000000000100","000000000000011101","000000000000010111","000000000000101010","000000000000100100","000000000000001000","111111111111100100","000000000000001011","111111111111110101","000000000000011101","000000000000100100","000000000000010000","000000000000001010","111111111111110111","000000000000010000","000000000000011001","111111111111010100","000000000000000100","111111111111101101","000000000000001100","111111111111101011","000000000000011110","111111111111110110","111111111111000101","111111111111111010","000000000000110100","111111111111110100","111111111111111101","111111111111110110","111111111111110001","000000000000110111","111111111111100101","000000000000001010","000000000000001110","000000000000001100","000000000000000111","000000000000001000","000000000000000101","000000000000010101","000000000000000111","000000000000000011","111111111111001111","111111111111110111","000000000000100110","000000000000100101","000000000000001011","111111111111101110","000000000000000000","111111111111111101","111111111111011001","111111111111110001","000000000000100000","000000000000000000","000000000000000001","111111111111100011","000000000000000000","111111111111100110","111111111111111010","111111111111001001","111111111111111100","111111111111101001","000000000000000000","111111111111011011","000000000000010100","000000000000000000","111111111111101011","111111111111010101","000000000000000101","111111111111101000","000000000000001000","000000000000100000","111111111111111101","000000000000001110","111111111111101010","000000000000010111","000000000000001011","000000000000011100","000000000000011100","111111111111101011","111111111111011011","000000000000100001","000000000000101110","111111111111010001","111111111111000110","000000000000010000","111111111111101010","111111111111111001","000000000000001010","000000000000010000","000000000000000010","111111111111100110","111111111111111001","111111111111101100","111111111111010110","111111111111111010","111111111111101011","000000000000000010","000000000000011100","111111111111101010","111111111111010110","111111111111110011","000000000000000001","111111111111101101","000000000000001010","111111111111111010","000000000000010100","000000000000001111","111111111111111110","000000000000001010","111111111111110100","000000000000001101","000000000000011001","111111111111111100","000000000000000000","111111111111010011","000000000000000001","111111111111111001","000000000000000000","000000000000000111","111111111111110000","000000000000100100","000000000000000100","000000000000010101","000000000000100110","111111111111110111","000000000000001110","000000000000110000","000000000000000000"),
("111111111111101001","000000000000001000","000000000000000000","000000000000100100","000000000000010011","111111111111110001","111111111111101100","000000000000010000","000000000000000111","111111111111111011","000000000000101010","000000000000001010","000000000000000111","000000000000000001","000000000000001001","000000000000001011","111111111111101011","000000000000000111","000000000000011100","111111111111101000","000000000000000011","000000000000100101","111111111111100101","111111111111100111","000000000000001010","000000000000011001","000000000000000101","111111111111111100","111111111111100000","111111111111110010","000000000000011110","111111111111101100","111111111111111010","111111111111011100","000000000000010100","000000000000010001","000000000000001111","000000000000010011","000000000000001101","111111111111101011","000000000000000000","111111111111011001","111111111111111000","000000000000011111","000000000000010000","111111111111110111","000000000000000111","111111111111100110","111111111111110000","111111111111101111","111111111111010010","000000000000011011","000000000000001010","000000000000001011","111111111111110111","000000000000011110","111111111111110100","111111111111101001","111111111111101110","111111111111111101","111111111111011110","111111111111111001","111111111111001010","111111111111110111","111111111111101111","000000000000001000","111111111111010110","111111111111011111","111111111111110100","000000000000000111","000000000000000100","111111111111110011","111111111111111101","111111111111101001","000000000000011000","111111111111101111","000000000000100000","000000000000000111","111111111111110101","111111111111101001","000000000000000011","000000000000001001","111111111110111100","111111111111010110","111111111111111101","000000000000000100","000000000000010111","111111111111100001","000000000000000000","111111111111100011","000000000000001001","111111111111110101","000000000000011001","111111111111100100","000000000000010001","111111111111110000","000000000000001111","000000000000011010","000000000000001111","111111111111011010","000000000000000001","000000000000100101","111111111111110111","000000000000100011","000000000000001101","000000000000001110","000000000000010010","111111111111111100","111111111111100110","111111111111111110","000000000000001001","000000000000000111","000000000000001000","000000000000010011","111111111111100001","111111111111100011","111111111111101100","111111111111100000","111111111111101011","111111111111111001","000000000000010100","111111111111111010","000000000000001011","000000000000100111","111111111111011101","000000000000011110","000000000000100110","000000000000010001"),
("111111111111110000","000000000000100110","000000000000010011","000000000000001010","000000000000001101","111111111111111100","000000000000010010","000000000000110001","000000000000001101","000000000000000101","000000000000010010","000000000000000100","000000000000000101","000000000000001101","000000000000010011","000000000000001110","111111111111101001","111111111111110000","111111111111111001","111111111111100101","111111111111101011","000000000000010011","111111111111100100","111111111111110100","000000000000010010","000000000000101001","111111111111111101","000000000000001111","111111111111100101","111111111111111110","000000000000100001","000000000000000111","000000000000001011","111111111111101011","000000000000000010","000000000000001010","111111111111110000","111111111111111000","000000000000000100","111111111111101000","111111111111110000","111111111111110101","111111111111100101","000000000000000100","000000000000100100","000000000000001111","000000000000001010","111111111111101010","111111111111101010","111111111111110110","111111111111101100","000000000000000011","111111111111101000","000000000000001101","111111111111100101","000000000000010101","111111111111101101","111111111111111101","000000000000001001","111111111111110111","111111111111101110","000000000000000100","111111111111010011","111111111111101010","111111111111011011","000000000000011100","111111111111101000","111111111111101010","000000000000010110","111111111111101101","000000000000000110","111111111111110110","111111111111110101","111111111111100101","000000000000101000","111111111111110011","000000000000010110","000000000000011110","000000000000010010","111111111111110000","000000000000010001","000000000000011100","111111111111100001","111111111111011101","111111111111101110","000000000000011001","111111111111110010","111111111111101011","111111111111101101","111111111111100000","000000000000000010","111111111111111001","000000000000010100","111111111111010100","000000000000011000","111111111111100110","000000000000000101","000000000000110001","000000000000001001","111111111111111010","111111111111111110","111111111111111010","111111111111010100","000000000000010000","111111111111101111","111111111111100110","000000000000100011","111111111111111100","000000000000000011","111111111111111000","000000000000100110","000000000000010111","000000000000000000","111111111111101111","111111111111101111","111111111111100111","000000000000001000","111111111111101011","000000000000000000","111111111111110101","111111111111111100","111111111111110010","000000000000001100","000000000000001011","111111111111101110","000000000000010100","000000000000001011","000000000000101011"),
("111111111111111110","000000000000001011","000000000000010010","000000000000001011","000000000000100111","000000000000001010","111111111111101101","000000000000100010","000000000000011000","000000000000000000","000000000000000100","111111111111100111","000000000000010111","000000000000010110","000000000000000011","111111111111111010","111111111111111100","000000000000011010","111111111111110111","111111111111101011","111111111111011101","000000000000000101","111111111111100101","111111111111111010","111111111111100011","000000000000100110","000000000000000101","000000000000100000","111111111111101111","000000000000001011","000000000000001101","111111111111111001","000000000000000000","111111111111101111","111111111111110000","000000000000010110","111111111111111110","000000000000011011","111111111111101100","000000000000000001","000000000000010001","111111111111110111","000000000000010110","000000000000011111","000000000000011100","000000000000000101","000000000000001011","111111111111110011","000000000000000000","111111111111011011","111111111111101000","000000000000011000","111111111111110111","000000000000011011","000000000000010000","000000000000010100","111111111111100001","111111111111111000","111111111111101001","111111111111110001","111111111111100010","000000000000010011","000000000000000010","000000000000000100","000000000000001000","111111111111111011","111111111111011010","111111111111101101","000000000000010011","000000000000011110","000000000000100100","000000000000000101","111111111111100000","111111111111101111","111111111111110100","000000000000001100","000000000000001000","000000000000000101","000000000000001110","111111111111110010","000000000000000010","000000000000011010","111111111111101110","111111111111111110","000000000000000100","000000000000000100","111111111111111100","000000000000000001","111111111111101000","111111111111111100","111111111111110111","111111111111111001","111111111111110000","111111111111110100","000000000000000100","111111111111100010","111111111111010111","000000000000100011","000000000000010101","000000000000001110","111111111111111000","111111111111110111","111111111111100111","000000000000001010","000000000000001101","000000000000000010","000000000000000100","111111111111101011","111111111111111010","111111111111100100","000000000000011010","000000000000010001","000000000000000000","111111111111110010","000000000000010111","111111111111100110","111111111111111011","111111111111011100","111111111111110000","000000000000000011","000000000000000100","111111111111010110","111111111111110000","000000000000011111","111111111111111110","000000000000000001","000000000000000000","000000000000001010"),
("000000000000000101","000000000000001100","000000000000010111","000000000000001000","111111111111111100","000000000000001001","111111111111111000","000000000000010111","111111111111101100","111111111111101000","000000000000001101","111111111111110001","111111111111110011","000000000000011010","111111111111101011","111111111111111011","111111111111110111","111111111111110011","111111111111110000","111111111111101110","111111111111011110","111111111111101111","111111111111100111","000000000000000111","000000000000001101","000000000000110000","000000000000011011","000000000000010110","111111111111110010","111111111111111111","000000000000011010","111111111111111001","000000000000100110","111111111111110011","111111111111110000","000000000000000011","111111111111111011","111111111111111110","000000000000000000","111111111111110000","111111111111100101","111111111111111000","111111111111101100","000000000000000000","000000000000111010","000000000000000001","111111111111011010","111111111111011000","111111111111101011","111111111111101101","111111111111100111","000000000000001000","111111111111100010","000000000000011100","000000000000000101","000000000000001110","111111111111110001","111111111111011101","111111111111110100","111111111111111001","111111111111011101","111111111111111011","111111111111101101","000000000000000000","000000000000011001","111111111111111100","111111111111101111","111111111111101010","000000000000000000","111111111111110101","000000000000011001","111111111111100111","111111111111010001","000000000000001101","000000000000000011","111111111111110111","000000000000100010","000000000000001110","000000000000001110","000000000000000011","000000000000011011","000000000000100100","111111111111010001","111111111111101111","111111111111110111","000000000000001111","111111111111111101","000000000000011010","111111111111111101","111111111111110111","111111111111111000","000000000000000110","111111111111111100","000000000000000000","111111111111111110","111111111111110001","111111111111011011","000000000000010110","000000000000100001","000000000000010011","111111111111110110","111111111111111100","111111111111111011","000000000000010101","111111111111110000","111111111111111100","000000000000000010","111111111111110101","111111111111111100","000000000000000101","000000000000011001","000000000000001111","111111111111110101","111111111111111000","000000000000001000","111111111111110001","111111111111111010","111111111111001111","000000000000001001","111111111111100011","111111111111110101","000000000000000101","111111111111110111","000000000000010100","111111111111100010","111111111111110111","000000000000000000","000000000000000100"),
("000000000000100000","000000000000100010","000000000000100100","000000000000011000","111111111111110000","000000000000000000","111111111111111001","000000000000011100","111111111111111010","111111111111011010","000000000000011111","111111111111110011","000000000000000101","000000000000100100","111111111111101001","000000000000001011","111111111111101101","111111111111111101","111111111111110111","111111111111110001","000000000000001001","111111111111111010","111111111111110110","000000000000011001","000000000000011011","000000000000001000","111111111111110000","000000000000010000","111111111111101101","111111111111110100","000000000000011011","111111111111100101","000000000000100001","111111111111100100","111111111111111011","111111111111111110","111111111111110001","000000000000000000","000000000000010000","111111111111100100","000000000000000001","111111111111101111","000000000000000011","000000000000010001","000000000000100101","111111111111111111","111111111111001011","111111111111110101","111111111111101001","000000000000000010","111111111111100101","000000000000000101","111111111111011001","000000000000101100","111111111111111011","111111111111110111","000000000000010101","111111111111101101","000000000000001000","000000000000010000","111111111111101000","000000000000010001","111111111111110100","000000000000000011","000000000000100011","000000000000001001","111111111111100011","000000000000000000","000000000000001110","111111111111111010","000000000000100011","111111111111010011","111111111111011010","111111111111110011","111111111111110111","000000000000000001","000000000000101001","000000000000011111","000000000000000000","111111111111010010","000000000000101000","000000000000110010","111111111111111001","111111111111100011","000000000000011000","111111111111111111","000000000000010111","111111111111111000","111111111111111110","111111111111100100","000000000000001111","000000000000010010","000000000000001100","111111111111100101","000000000000001011","000000000000011010","111111111111011111","000000000000111010","000000000000100010","111111111111110011","000000000000010000","111111111111101100","111111111111100100","111111111111110000","111111111111110100","111111111111100111","000000000000010011","111111111111001110","000000000000000000","111111111111100100","000000000000001001","000000000000110111","000000000000001101","111111111111000111","111111111111111011","111111111111111111","000000000000000100","111111111111100010","000000000000100110","111111111111110010","111111111111100010","000000000000000001","000000000000010010","000000000000000000","111111111111001010","000000000000001010","111111111111100001","000000000000010001"),
("000000000000010101","111111111111110011","111111111111110111","000000000000000101","000000000000000000","000000000000001101","000000000000011011","111111111111110000","111111111111110110","000000000000001010","000000000000001111","111111111111101010","000000000000010100","000000000000010100","111111111111011001","000000000000100011","111111111111110010","000000000000011111","111111111111110000","000000000000001000","000000000000000011","000000000000000010","000000000000011010","111111111111111110","000000000000000111","000000000000000001","111111111111111100","000000000000111110","000000000000001000","111111111111111001","000000000000011011","111111111111101100","000000000000011011","111111111111110010","111111111111111110","111111111111010101","000000000000011000","000000000000010000","111111111111101010","000000000000000111","000000000000001101","111111111111110001","000000000000010101","000000000000000101","111111111111101011","111111111111110110","111111111111100000","111111111111101100","111111111111100001","111111111111110100","000000000000000111","000000000000000011","111111111111111111","000000000000010100","000000000000001010","111111111111101100","111111111111111000","000000000000000111","111111111111111001","000000000000010001","111111111111110110","000000000000001101","111111111111111001","111111111111101000","000000000000011011","111111111111101110","111111111111011100","000000000000000110","000000000000010011","111111111111110011","000000000000011000","111111111111101111","111111111111101001","000000000000000010","000000000000001000","000000000000100100","000000000000010111","000000000000011010","000000000000000101","111111111111100000","111111111111111000","000000000000000111","111111111111111100","111111111111001011","000000000000100100","111111111111101101","000000000000001010","000000000000001110","111111111111101010","111111111111100011","111111111111110100","000000000000010010","000000000000000011","000000000000000000","111111111111101100","000000000000001101","111111111111110110","000000000000110010","000000000000000011","111111111111111010","000000000000010101","111111111111010001","111111111111110101","111111111111101100","111111111111100110","111111111111101100","111111111111111000","111111111111100000","111111111111010111","111111111111110010","000000000000000000","000000000000110010","111111111111100010","111111111111011010","111111111111011010","111111111111110011","111111111111110011","000000000000010001","111111111111110111","000000000000000110","000000000000011111","000000000000010011","000000000000001100","000000000000110011","111111111111100000","000000000000001010","000000000000100000","111111111111101100"),
("111111111111111100","111111111111101000","111111111111110110","000000000000001111","111111111111111000","000000000000000111","000000000000000000","000000000000010001","000000000000000110","000000000000001001","000000000000001111","111111111111101100","000000000000011111","111111111111111111","000000000000000000","000000000000011011","000000000000011001","111111111111111100","111111111111101110","000000000000000111","111111111111100100","111111111111110011","111111111111111110","111111111111110110","111111111111111001","000000000000001100","111111111111110011","000000000000000000","111111111111110100","000000000000100001","000000000000001000","111111111111110010","000000000000010110","111111111111011101","000000000000000111","000000000000010001","000000000000000000","111111111111111011","000000000000000110","000000000000000010","111111111111011010","111111111111110100","000000000000010011","000000000000001110","000000000000010010","111111111111110101","111111111111111011","111111111111111100","111111111111011000","111111111111111000","111111111111101111","000000000000001010","111111111111101000","111111111111110101","000000000000100010","000000000000011100","111111111111111011","000000000000001100","111111111111111110","000000000000000100","111111111111100000","000000000000010100","000000000000010110","000000000000010100","111111111111101000","111111111111111100","111111111111101000","000000000000000111","000000000000001111","111111111111110010","111111111111111111","000000000000001000","111111111111101100","000000000000000111","111111111111100110","000000000000000110","000000000000000111","000000000000000011","000000000000000000","111111111111111101","111111111111110110","000000000000000100","000000000000010000","111111111111111000","111111111111111111","000000000000001001","000000000000000101","000000000000010111","111111111111111100","000000000000001000","000000000000001100","111111111111111010","111111111111101011","000000000000010100","111111111111111111","111111111111111001","111111111111110000","000000000000000000","000000000000010100","000000000000000000","000000000000010111","111111111111111100","111111111111110010","111111111111110010","111111111111111100","000000000000001011","111111111111110110","111111111111100000","111111111111101010","111111111111111000","111111111111100101","000000000000000110","000000000000001011","111111111111110111","000000000000000001","111111111111101000","111111111111110100","111111111111100001","111111111111110000","000000000000000011","000000000000000011","000000000000000110","000000000000100000","000000000000001000","000000000000000000","111111111111110001","000000000000011100","111111111111110000"),
("000000000000000000","000000000000000010","111111111111101010","111111111111111111","000000000000010000","111111111111111111","111111111111111111","000000000000000010","000000000000010001","111111111111110111","000000000000010100","111111111111010101","000000000000000001","111111111111110010","000000000000001010","000000000000001111","000000000000001011","000000000000010100","111111111111110100","000000000000010111","000000000000001000","000000000000001111","000000000000010100","111111111111101111","111111111111110110","111111111111111000","000000000000001111","111111111111111101","000000000000001110","000000000000010010","000000000000010011","111111111111110000","111111111111110001","000000000000010011","111111111111111101","000000000000001110","000000000000000010","000000000000001111","000000000000000001","111111111111100111","111111111111111100","111111111111101111","111111111111111001","000000000000010100","111111111111111100","000000000000011010","000000000000010100","000000000000000110","111111111111100000","111111111111111111","111111111111110001","000000000000000100","000000000000000101","111111111111111011","111111111111111011","000000000000010101","111111111111111010","111111111111110011","111111111111111111","000000000000000111","000000000000000011","111111111111111101","000000000000001111","111111111111101000","000000000000000000","000000000000000111","111111111111101001","111111111111111001","111111111111110101","111111111111111101","000000000000000001","000000000000011001","000000000000010101","000000000000000000","111111111111101010","000000000000010010","000000000000000110","111111111111110111","111111111111110110","000000000000001101","111111111111111101","111111111111100101","000000000000011100","000000000000010000","000000000000001110","000000000000001101","000000000000010011","000000000000010010","000000000000000100","000000000000100001","000000000000000111","111111111111110011","111111111111101100","000000000000000011","111111111111111001","111111111111110100","111111111111101110","111111111111111111","000000000000001011","000000000000001111","111111111111111011","111111111111111111","111111111111101010","000000000000011000","000000000000010101","000000000000001001","111111111111110101","000000000000001011","000000000000000000","000000000000000010","111111111111110101","000000000000010000","000000000000000000","111111111111111110","111111111111111011","111111111111111111","111111111111111000","000000000000011111","000000000000000111","000000000000010001","111111111111111011","000000000000011000","000000000000011100","000000000000001101","000000000000010100","111111111111110010","111111111111111000","000000000000000101"),
("000000000000000111","111111111111111100","000000000000010001","111111111111110101","111111111111101101","000000000000001000","000000000000010100","000000000000001100","111111111111111111","000000000000001000","000000000000000000","000000000000001001","111111111111110011","111111111111111111","000000000000001001","000000000000001000","111111111111101110","000000000000001001","000000000000001010","000000000000001101","111111111111111000","111111111111110111","000000000000010000","000000000000001001","111111111111111101","000000000000000011","000000000000001100","000000000000000110","000000000000001100","111111111111111011","000000000000001110","111111111111101101","111111111111110001","000000000000001011","000000000000000110","111111111111111010","111111111111110001","111111111111111100","000000000000001000","111111111111111000","111111111111111000","000000000000010010","000000000000010010","000000000000010011","111111111111111000","000000000000001010","111111111111111001","111111111111110110","000000000000010001","111111111111110111","111111111111111101","111111111111110110","111111111111101111","000000000000001111","000000000000000001","000000000000000000","000000000000010011","111111111111111010","111111111111111111","000000000000010001","111111111111110000","000000000000010000","111111111111111100","000000000000001100","000000000000000000","000000000000000000","111111111111101110","111111111111110011","111111111111111001","111111111111110111","111111111111101101","111111111111111101","111111111111111101","000000000000001101","111111111111111001","111111111111101110","000000000000001001","111111111111110011","000000000000010000","000000000000000011","111111111111110011","000000000000001001","000000000000000110","000000000000001111","111111111111101100","111111111111110001","111111111111111010","111111111111101111","000000000000001100","111111111111110011","111111111111111011","000000000000001011","000000000000000010","000000000000001110","111111111111110110","111111111111101100","111111111111110111","000000000000010011","111111111111110001","000000000000001011","111111111111110111","000000000000000111","111111111111111111","111111111111101110","111111111111101100","111111111111110001","000000000000000010","000000000000001100","111111111111101101","111111111111111101","111111111111110110","111111111111111100","111111111111111000","111111111111110100","111111111111101101","111111111111101100","111111111111101110","000000000000000111","000000000000001100","111111111111110000","111111111111111110","111111111111111001","000000000000001111","000000000000001010","000000000000000110","000000000000001111","000000000000001111","111111111111111100"),
("111111111111110111","111111111111110110","000000000000000011","111111111111110000","000000000000000010","111111111111101101","111111111111110000","000000000000010010","000000000000000110","111111111111111100","000000000000010100","000000000000000101","111111111111101100","111111111111110100","111111111111101101","111111111111101100","111111111111110110","000000000000001011","111111111111110001","111111111111110001","111111111111111111","000000000000000000","111111111111111001","000000000000001111","000000000000001111","000000000000000110","111111111111101110","000000000000010000","111111111111110001","111111111111111000","000000000000010010","111111111111111101","111111111111111100","000000000000001100","111111111111111000","111111111111101100","111111111111110100","111111111111111010","000000000000010001","111111111111111010","000000000000001000","111111111111111100","000000000000001111","000000000000000000","000000000000001000","111111111111111101","000000000000001011","000000000000001100","000000000000010001","000000000000000101","000000000000000011","111111111111111010","000000000000001111","000000000000000001","000000000000000101","000000000000000010","111111111111101101","000000000000001110","000000000000010100","111111111111111101","111111111111111101","000000000000001110","111111111111110000","111111111111110001","000000000000000101","111111111111111010","111111111111110001","000000000000001111","000000000000000000","111111111111110110","111111111111110110","000000000000010100","000000000000001011","000000000000001010","000000000000001000","111111111111111100","000000000000001101","000000000000000100","111111111111110010","000000000000001111","111111111111110000","000000000000000011","000000000000000010","000000000000000010","111111111111111010","000000000000001000","111111111111111000","000000000000000001","000000000000000000","000000000000000010","111111111111111111","000000000000010010","111111111111111101","000000000000001001","111111111111101111","111111111111111010","111111111111101110","111111111111111000","111111111111111011","000000000000000000","000000000000010001","111111111111101100","000000000000000001","111111111111110000","111111111111110101","000000000000001111","000000000000000010","000000000000010100","111111111111111011","111111111111110000","000000000000010100","111111111111101110","111111111111110110","000000000000010010","111111111111110111","000000000000001100","000000000000001001","111111111111101101","000000000000001001","111111111111111110","111111111111111000","000000000000000011","111111111111111101","111111111111111001","000000000000000110","111111111111111010","111111111111101100","111111111111101110"),
("111111111111111001","000000000000001111","111111111111111101","000000000000000010","111111111111101111","111111111111111110","000000000000010011","000000000000001001","000000000000010100","111111111111110011","111111111111111110","000000000000000010","111111111111101111","111111111111101111","000000000000001010","111111111111110111","111111111111110011","000000000000000100","111111111111110110","000000000000010010","111111111111110011","000000000000010011","111111111111111110","111111111111111000","000000000000001001","000000000000000110","000000000000010100","111111111111111111","000000000000001111","000000000000010011","000000000000000010","111111111111111010","000000000000000000","000000000000010000","111111111111111000","000000000000010100","000000000000000010","000000000000010001","111111111111110010","000000000000000111","000000000000000100","111111111111111110","000000000000010100","111111111111101110","000000000000000000","111111111111101110","000000000000010001","000000000000001101","000000000000010011","111111111111110100","000000000000001100","111111111111110010","111111111111111110","111111111111111000","111111111111111111","111111111111110001","111111111111101101","000000000000010000","000000000000010001","000000000000001100","111111111111110110","000000000000000000","111111111111110001","000000000000000001","111111111111110101","000000000000001010","111111111111101101","000000000000000100","111111111111110010","111111111111111000","000000000000001110","000000000000000100","111111111111101110","111111111111111100","111111111111111001","000000000000010010","000000000000000000","111111111111110011","111111111111110010","111111111111111101","111111111111101111","000000000000010001","111111111111111111","111111111111110010","000000000000000011","111111111111110101","000000000000001000","000000000000010100","000000000000000110","000000000000000010","111111111111111101","111111111111111111","000000000000001011","111111111111111111","000000000000001011","000000000000000010","111111111111101111","111111111111111111","111111111111111010","111111111111110000","111111111111101110","111111111111110000","000000000000001111","111111111111110111","000000000000000101","000000000000000001","000000000000001001","111111111111111110","000000000000000010","000000000000000011","000000000000000000","000000000000010001","111111111111110111","000000000000000011","111111111111110101","111111111111110011","000000000000001100","000000000000000110","111111111111101111","111111111111111001","000000000000001100","000000000000010001","000000000000000011","000000000000000110","000000000000010100","111111111111111010","000000000000001000","000000000000000010"),
("000000000000010100","000000000000000011","000000000000000010","000000000000010011","111111111111100100","000000000000010010","111111111111101110","000000000000001000","111111111111111000","000000000000000110","111111111111101111","000000000000001000","000000000000000010","000000000000010111","111111111111100011","111111111111110001","000000000000001101","111111111111011000","111111111111111000","000000000000001010","111111111111101110","111111111111101001","111111111111101010","000000000000010000","111111111111111100","000000000000001111","111111111111101001","000000000000101001","111111111111101011","111111111111110000","111111111111111111","000000000000011011","000000000000001011","000000000000000011","111111111111111101","000000000000001000","111111111111100000","000000000000001110","000000000000010000","111111111111101011","111111111111100110","000000000000000000","000000000000000011","000000000000000100","000000000000011111","000000000000000010","000000000000000011","111111111111010100","111111111111011010","000000000000001010","111111111111110111","000000000000010100","000000000000000000","000000000000010010","111111111111111100","111111111111101110","000000000000001010","000000000000001011","000000000000000011","000000000000001100","000000000000100111","000000000000010110","111111111111101010","111111111111111111","000000000000000110","111111111111110101","000000000000001011","000000000000001011","111111111111111111","111111111111110001","000000000000001000","000000000000001000","000000000000001110","000000000000000001","000000000000000000","000000000000010111","111111111111101111","000000000000001011","111111111111011101","111111111111111010","000000000000001101","000000000000000000","000000000000001101","111111111111100000","000000000000100001","111111111111101110","111111111111011101","000000000000000100","000000000000000111","000000000000010011","111111111111110010","000000000000100101","000000000000000011","111111111111111110","111111111111101000","000000000000001101","000000000000010001","000000000000010011","000000000000000101","111111111111110100","000000000000000111","000000000000001000","000000000000000011","000000000000010010","111111111111100100","111111111111110000","000000000000000010","111111111111111011","111111111111111101","111111111111111010","000000000000001000","000000000000010111","000000000000000110","111111111111101000","000000000000001011","000000000000000110","000000000000010011","000000000000000001","000000000000010101","000000000000011111","111111111111101111","111111111111110110","000000000000001001","111111111111111010","111111111111111111","000000000000010100","111111111111010011","000000000000001101"),
("000000000000100101","111111111111101110","000000000000100111","111111111111101011","000000000000000010","111111111111110100","000000000000010111","111111111111111111","111111111111101100","111111111111101010","111111111111011000","000000000000010010","000000000000000111","000000000000000110","111111111111111011","000000000000000101","000000000000010011","111111111111111011","000000000000010111","000000000000000100","000000000000010010","000000000000011100","000000000000011001","111111111111111101","000000000000000101","111111111111110100","000000000000000010","111111111111101000","000000000000000000","000000000000011010","000000000000001010","111111111111110101","111111111111100111","000000000000000010","000000000000001111","111111111111101001","000000000000000011","111111111111100110","000000000000011001","000000000000000000","000000000000100100","000000000000000100","000000000000001011","111111111111101111","111111111111101100","000000000000000000","000000000000010101","000000000000001110","000000000000001000","000000000000000011","111111111111111110","111111111111110010","000000000000001001","111111111111111101","000000000000010000","111111111111110110","000000000000100010","111111111111111101","000000000000010000","000000000000000010","111111111111110111","000000000000011001","000000000000011000","111111111111101101","000000000000000000","000000000000001111","000000000000000000","111111111111111011","000000000000000110","000000000000010011","111111111111101000","111111111111111000","111111111111111111","111111111111100111","111111111111110110","111111111111110011","000000000000010101","111111111111011100","000000000000001111","111111111111110100","111111111111111111","111111111111110011","111111111111110001","000000000000000110","111111111111111101","000000000000010100","000000000000010000","111111111111110100","111111111111011110","000000000000010101","111111111111111000","111111111111111001","000000000000010010","111111111111111011","000000000000000000","111111111111101011","000000000000000000","000000000000001110","000000000000001110","000000000000001000","111111111111101000","000000000000100011","111111111111111100","111111111111100101","000000000000010101","111111111111101111","000000000000000000","000000000000000001","000000000000000101","000000000000001111","000000000000000000","000000000000001001","000000000000000000","000000000000001000","111111111111111000","111111111111101010","111111111111100110","000000000000001000","111111111111101111","111111111111110001","000000000000010001","111111111111111010","111111111111111011","111111111111011000","000000000000011110","000000000000001011","000000000000101011","111111111111110000"),
("111111111111100001","111111111111101101","000000000000001111","111111111111010100","111111111111011111","111111111111101011","000000000000000100","111111111111111101","111111111111101101","000000000000001110","111111111111110001","111111111111111010","000000000000000101","000000000000110000","111111111111101111","111111111111100100","000000000000001110","111111111111101110","000000000000000011","000000000000101000","111111111111111000","000000000000100111","000000000000100111","111111111111100100","000000000000010100","111111111111110010","111111111111110110","111111111111101000","000000000000001001","000000000000001010","111111111111110011","000000000000100101","000000000000010100","000000000000010100","000000000000001110","111111111111101010","000000000000010111","111111111111011101","000000000000000001","000000000000100010","000000000000010011","111111111111111011","000000000000001101","111111111111011000","000000000000000111","111111111111111001","111111111111100010","111111111111110010","000000000000010100","000000000000011011","111111111111100010","111111111111100001","111111111111111101","000000000000010000","000000000000110001","000000000000000111","000000000000011010","000000000000011111","111111111111111100","111111111111111011","000000000000001101","000000000000010010","111111111111111100","111111111111010000","000000000000000110","000000000000000000","111111111111100001","111111111111101101","000000000000011111","000000000000000111","111111111111101101","111111111111101010","000000000000011101","000000000000001000","111111111111110111","000000000000010011","111111111111100010","000000000000010001","000000000000010101","000000000000001110","111111111111100010","111111111111110000","111111111111111100","000000000000101000","111111111111010010","000000000000010111","000000000000000011","000000000000010110","000000000000000110","000000000000010101","000000000000000110","111111111111110011","000000000000000111","000000000000100010","000000000000000000","111111111111111110","000000000000011010","000000000000111001","000000000000000111","000000000000001100","111111111111100110","000000000000000000","000000000000001000","111111111111010110","000000000000000011","111111111111001110","000000000000001000","000000000000010110","000000000000100010","000000000000010110","000000000000000011","111111111111111110","111111111111010111","000000000000000010","111111111111101100","111111111111111110","111111111111110000","000000000000100101","111111111111111010","111111111111111111","000000000000001110","111111111111101010","000000000000010110","111111111111101001","000000000000011011","111111111111110111","111111111111111010","000000000000001101"),
("111111111111111000","111111111111101011","000000000000011010","111111111111100110","111111111111011111","111111111111111010","000000000000001011","111111111111010110","000000000000010001","111111111111110011","111111111111101011","111111111111110101","111111111111101100","000000000000010100","111111111111010100","111111111110111111","111111111111100110","111111111111001110","111111111111011011","000000000000000110","111111111111100001","000000000000101101","000000000000000010","111111111111010001","000000000000000000","111111111111100101","111111111111001110","111111111111110001","000000000000010000","000000000000000001","111111111111101011","000000000000011001","000000000000100110","111111111111111000","111111111111110100","111111111111011010","000000000000001000","111111111111101010","000000000000101111","000000000000010111","111111111111101000","111111111111110100","000000000000101100","111111111111100111","111111111111110101","000000000000010101","111111111111100001","111111111111101111","111111111111110110","000000000000110111","111111111111100110","111111111111101100","111111111111110011","000000000000011111","000000000000101001","000000000000011010","000000000000011101","000000000000001110","000000000000010000","000000000000010010","000000000000010111","000000000000011000","000000000000000011","111111111111001111","111111111111101011","111111111111101101","111111111111100111","111111111111110000","000000000000110010","000000000000000010","000000000000000101","111111111111101110","000000000000110001","000000000000011101","000000000000100100","000000000000110110","111111111111111101","000000000000011000","000000000000001001","111111111111110011","111111111111110011","000000000000001101","000000000000011010","000000000000001000","111111111111011111","000000000000100100","111111111111110000","000000000000011000","000000000000001000","000000000000010110","000000000000000001","000000000000010111","000000000000000110","000000000000010110","000000000000010011","000000000000010001","000000000000100100","000000000000100011","111111111111110011","000000000000100001","111111111111110100","000000000000000110","000000000000011110","111111111111010000","111111111111001010","111111111111010001","000000000000010001","111111111111111110","000000000000111001","000000000000010010","111111111111110111","111111111111101111","111111111111011110","000000000000001100","000000000000100001","111111111111111110","000000000000000000","000000000000000100","000000000000000101","000000000000001111","000000000000000101","111111111111101101","111111111111101101","111111111111010111","000000000000010111","111111111111100101","111111111111101110","000000000001000100"),
("111111111111111010","111111111111101111","000000000000001100","000000000000000100","111111111111010000","111111111111111000","111111111111111101","111111111111001000","000000000000101110","000000000000001011","111111111111111101","000000000000010000","000000000000000011","000000000000000100","111111111111100110","111111111111010100","111111111111101000","111111111111101100","111111111111111001","000000000000100111","111111111111011010","000000000000011010","111111111111011100","111111111111110111","111111111111110001","111111111111110101","111111111111001011","000000000000001000","000000000000100000","111111111111111110","111111111111111011","000000000000101001","000000000000100111","000000000000000011","111111111111110000","111111111111100011","111111111111111010","000000000000010011","111111111111101101","111111111111111001","111111111111100010","111111111111111110","111111111111110101","111111111110111100","000000000000011010","000000000000100011","000000000000001010","111111111111100000","000000000000010100","000000000000101110","111111111111010110","000000000000000110","111111111111111111","000000000000000111","000000000000101010","111111111111111000","111111111111111001","000000000000011001","111111111111111001","000000000000010000","000000000000101011","000000000000001101","111111111111101000","111111111111101000","111111111111011100","111111111111100100","111111111111000000","111111111111111110","000000000000101011","111111111111110110","000000000000001100","000000000000011000","000000000000010001","111111111111111001","000000000000110111","000000000000001110","000000000000000100","000000000000000000","000000000000010000","111111111111111010","111111111111110000","000000000000000000","111111111111111001","111111111111001111","000000000000001100","111111111111101011","000000000000000101","000000000000000111","000000000000010101","000000000000011000","111111111111101100","000000000000011001","111111111111111010","111111111111101110","111111111111111010","000000000000010010","000000000000101001","000000000000100100","111111111111111001","000000000000011111","000000000000000001","000000000000000000","000000000000101000","111111111111111101","111111111111110110","111111111111101010","000000000000001010","000000000000000001","000000000000010111","111111111111101000","111111111111110100","111111111111110010","111111111111111001","000000000000101110","000000000000010010","000000000000011100","000000000000001000","000000000000010111","111111111111101001","000000000000010010","000000000000001000","111111111111110101","111111111111100101","000000000000000101","000000000000001000","000000000000001101","111111111111101001","000000000000100110"),
("000000000000001001","111111111111110100","000000000000000101","111111111111110110","111111111111011000","111111111111101100","111111111111101111","111111111111001010","000000000000101011","000000000000001010","000000000000000001","000000000000100001","000000000000001100","000000000000000000","111111111111011000","111111111111100010","111111111111001000","111111111111100111","000000000000011110","000000000000010111","111111111111110100","000000000000010101","111111111111101100","111111111111101010","000000000000000010","111111111111110011","111111111111000000","000000000000010011","000000000000010010","000000000000000100","111111111111111000","000000000000010101","000000000000011001","000000000000001010","111111111111101110","000000000000000000","111111111111101010","111111111111110010","111111111111110100","000000000000000110","000000000000001110","000000000000000101","111111111111010011","111111111111001111","111111111111111101","111111111111111100","111111111111001101","111111111111011101","000000000000000011","000000000000010011","111111111111011100","111111111111111011","000000000000000100","000000000000010100","000000000000011001","000000000000001110","111111111111111010","000000000000101110","000000000000000001","000000000000001001","000000000000100001","000000000000000000","111111111111111100","111111111111101111","111111111111101010","111111111111111010","111111111111100001","000000000000000001","000000000000111101","000000000000000101","111111111111111100","000000000000010000","000000000000010000","000000000000011001","000000000000100111","000000000000001000","111111111111110010","111111111111111111","000000000000000001","111111111111110011","111111111111101011","111111111111111110","111111111111111001","111111111111101101","000000000000010000","111111111111111000","000000000000010101","000000000000010010","000000000000001011","000000000000101000","111111111111011110","000000000000001000","111111111111011100","111111111111111010","000000000000000100","000000000000011010","000000000000000111","000000000000110101","111111111111101011","000000000000000011","111111111111101111","111111111111100001","000000000000100000","111111111111100100","111111111111111100","111111111111100110","000000000000001000","000000000000100010","000000000000010100","111111111111010111","000000000000011001","111111111111100110","000000000000010001","000000000000000110","000000000000010001","111111111111111110","000000000000010110","000000000000011001","111111111111101100","000000000000100110","000000000000011000","111111111111110110","000000000000010000","111111111111111011","111111111111110000","111111111111101100","111111111111111111","000000000000000110"),
("111111111111111110","000000000000001111","111111111111110101","000000000000010011","111111111111110111","111111111111101101","111111111111110110","111111111111100000","000000000000110001","111111111111111101","111111111111111011","000000000000011110","111111111111101010","000000000000001101","111111111111110100","111111111111100100","111111111111101111","111111111111100101","000000000000010101","000000000000011101","111111111111111000","000000000000000010","000000000000000111","111111111111101010","111111111111100100","111111111111110000","111111111111001110","000000000000100000","000000000000001101","000000000000001010","111111111111100011","000000000000101100","000000000000011101","000000000000000001","111111111111010101","000000000000000111","111111111111111100","111111111111110011","111111111111111000","000000000000010111","000000000000100100","111111111111111111","111111111111001100","111111111111011010","111111111111111001","000000000000000100","111111111111010001","111111111111010111","000000000000001101","000000000000101010","111111111111100010","111111111111110100","000000000000001110","000000000000010111","000000000000011100","111111111111111011","000000000000010110","000000000000101101","000000000000000010","111111111111110001","000000000000011000","000000000000101011","000000000000000000","111111111111110101","000000000000000101","111111111111011101","111111111111110000","111111111111101100","000000000001010110","111111111111101100","000000000000010000","000000000000010101","111111111111111001","000000000000010010","000000000000111110","000000000000001011","111111111111100010","000000000000010001","111111111111111010","111111111111100110","111111111111110101","111111111111110001","000000000000001001","111111111111111011","111111111111110111","111111111111111011","000000000000001001","000000000000011100","111111111111111100","000000000000010100","111111111111011111","000000000000100111","111111111111010000","111111111111110111","111111111111110111","000000000000000010","000000000000000010","000000000000011110","111111111111011100","000000000000010110","111111111111101110","111111111111110001","000000000000001000","111111111111101101","111111111111011100","111111111111011111","000000000000011110","000000000000000010","000000000000010001","111111111111011101","000000000000011011","111111111111011010","111111111111101010","000000000000000101","000000000000101001","000000000000010100","000000000000010110","000000000000101000","000000000000000101","000000000000110011","000000000000100110","111111111111010011","000000000000001110","000000000000001110","111111111111010010","111111111111110111","000000000000010001","000000000000010101"),
("111111111111111000","000000000000001100","000000000000010010","111111111111111110","111111111111010001","111111111111101001","111111111111110110","111111111111011001","111111111111111101","000000000000000011","111111111111101100","000000000000011010","111111111111010110","000000000000001000","111111111111110011","111111111111110011","111111111111100100","000000000000000111","000000000000001011","000000000000000011","111111111111110110","111111111111100010","111111111111110000","111111111111110101","000000000000000010","111111111111110011","111111111111101000","000000000000000011","000000000000000011","111111111111110101","111111111111101011","000000000000011001","000000000000001111","111111111111111110","111111111111110011","111111111111110010","000000000000000000","000000000000000101","000000000000010001","000000000000011010","000000000000101000","000000000000010011","111111111110100100","111111111111010011","000000000000010101","000000000000011111","111111111111111011","111111111111100101","000000000000011111","000000000000101011","111111111111111011","111111111111100001","000000000000011011","111111111111111111","000000000000000001","000000000000011000","000000000000110000","000000000000100000","000000000000010101","111111111111111010","000000000000101111","000000000000010010","000000000000000111","000000000000000101","000000000000000000","111111111111101101","111111111111110010","111111111111110000","000000000000110100","111111111111110101","111111111111111101","000000000000011011","111111111111100110","000000000000001000","000000000000011011","000000000000001000","111111111111100001","000000000000010100","000000000000000101","111111111111100101","111111111111100001","000000000000000110","111111111111010010","111111111111111000","111111111111110111","111111111111110100","111111111111101101","000000000000001111","000000000000010110","000000000000011100","111111111111111111","000000000000010110","111111111111100010","111111111111100001","111111111111110111","000000000000000111","000000000000001011","000000000000101001","000000000000010011","000000000000101100","111111111111111111","111111111111011110","000000000000100110","111111111111111000","000000000000000000","111111111111011111","000000000000010111","111111111111111010","000000000000011011","111111111111100010","000000000000100001","111111111111110101","000000000000001110","000000000000011100","000000000000001010","000000000000000001","000000000000000111","000000000000011110","111111111111110111","000000000000101011","000000000000011111","111111111111011011","111111111111110111","111111111111111110","111111111111101110","000000000000000110","000000000000011011","000000000000100110"),
("000000000000001000","000000000000011101","000000000000001010","111111111111111000","111111111110101000","111111111111101001","000000000000101010","111111111111010010","000000000000011000","111111111111111000","111111111111011011","000000000000100111","111111111111010101","111111111111110000","111111111111101101","111111111111110101","111111111111100100","111111111111101001","000000000000010100","111111111111111110","111111111111111111","111111111111011010","111111111111001101","000000000000010010","111111111111111100","000000000000010101","111111111111100011","000000000000010000","111111111111110111","111111111111111011","111111111111100001","111111111111111111","000000000000110000","000000000000000010","000000000000001001","000000000000000101","111111111111111101","000000000000000101","111111111111111110","000000000000001101","111111111111111001","000000000000000110","111111111110101100","111111111111010011","000000000000000110","000000000000001010","000000000000000000","111111111111101110","000000000000100011","000000000000101010","111111111111100011","111111111111110101","000000000000000101","000000000000100001","000000000000010100","000000000000000111","000000000000101001","000000000000101111","000000000000011101","111111111111101101","000000000000100001","000000000000011101","000000000000010100","000000000000000000","000000000000000000","000000000000011011","111111111111101010","111111111111111011","000000000000101110","111111111111111110","000000000000000101","000000000000001011","111111111111100100","000000000000000100","000000000000000010","000000000000001010","000000000000001101","000000000000010011","000000000000000111","111111111111110101","111111111111011000","000000000000001100","111111111111001111","000000000000000000","111111111111100111","111111111111110101","000000000000000011","111111111111101011","111111111111111100","000000000000010101","111111111111011111","000000000000000001","111111111111101010","111111111111000011","111111111111110111","000000000000000101","111111111111101111","000000000001010110","111111111111101111","000000000000101010","111111111111111100","111111111111101011","000000000000010011","111111111111101001","111111111111101011","111111111111100000","000000000000001000","000000000000110100","111111111111111010","111111111111110010","000000000000011100","111111111111100010","000000000000100100","000000000000101111","000000000000100100","000000000000000000","000000000000001001","000000000000000000","111111111111110011","000000000000100101","000000000000000110","000000000000000110","111111111111011111","111111111111001010","000000000000000111","111111111111110111","111111111111111110","000000000000001100"),
("000000000000000111","000000000000000101","000000000000101111","111111111111111110","111111111110111110","111111111111101101","000000000000001000","111111111111011101","111111111111110101","111111111111110011","111111111111001110","000000000000010111","111111111111110010","111111111111101101","000000000000001110","111111111111101001","111111111111011101","000000000000000011","000000000000011010","111111111111110100","111111111111110001","111111111111100100","111111111111000110","111111111111110001","000000000000011000","111111111111110010","111111111111111101","000000000000001110","111111111111110111","111111111111110010","000000000000000010","000000000000001111","000000000000110011","111111111111111101","111111111111111011","111111111111101001","000000000000010111","111111111111111011","000000000000000101","000000000000100011","000000000000001101","111111111111111011","111111111110101000","111111111111011000","111111111111111000","000000000000100010","111111111111100110","000000000000000100","000000000000101101","000000000000101011","111111111111111000","111111111111011111","000000000000000111","111111111111111000","111111111111111001","000000000000010110","000000000000100100","000000000000001100","000000000000100010","111111111111111110","000000000000011101","000000000000100110","000000000000001100","000000000000000011","111111111111011101","000000000000001100","111111111111011111","111111111111100111","000000000000011001","000000000000000000","000000000000001111","000000000000010001","111111111111110111","000000000000001101","000000000000011011","111111111111101101","111111111111101111","000000000000010011","000000000000000000","111111111111111001","111111111111110010","000000000000010101","000000000000001110","111111111111110011","111111111111011100","111111111111110100","000000000000000001","111111111111101110","111111111111101010","000000000000001001","000000000000000000","000000000000011001","111111111111100111","111111111111100101","000000000000001011","000000000000000100","111111111111101011","000000000001000000","111111111111100001","000000000000110100","111111111111111001","111111111111101111","000000000000011011","111111111111110011","000000000000010110","111111111111101101","000000000000010101","000000000000100011","111111111111100111","000000000000000000","000000000000010110","111111111111100100","111111111111110101","000000000000001100","000000000000101101","111111111111111110","000000000000010101","000000000000000111","000000000000000101","000000000000011111","000000000000001010","111111111111111001","111111111111111001","111111111111100101","000000000000000000","000000000000000010","000000000000100001","000000000000101011"),
("000000000000001011","111111111111111101","000000000000010010","000000000000011000","111111111111000100","111111111111101001","000000000000010001","000000000000001101","000000000000010011","000000000000001100","000000000000001011","000000000000011111","111111111111101100","111111111111101010","111111111111111010","111111111111111111","111111111111101101","111111111111101001","000000000000010100","111111111111111110","000000000000001111","111111111111010111","111111111110110010","111111111111101100","000000000000000111","000000000000011001","000000000000000101","000000000000100001","000000000000010000","111111111111111100","000000000000011000","000000000000011001","000000000000100001","111111111111110100","111111111111100100","111111111111111101","000000000000000111","111111111111111111","111111111111111001","000000000000100110","000000000000010110","111111111111111011","111111111111001001","111111111111100111","111111111111110101","000000000000011001","111111111111100101","111111111111100101","000000000000011011","000000000000010110","111111111111110000","111111111111101111","000000000000001101","000000000000000001","000000000000010110","111111111111110100","000000000000101001","000000000000011001","111111111111101110","000000000000001000","000000000000100111","000000000000011101","000000000000000001","111111111111111100","111111111111110001","111111111111101100","111111111111110011","111111111111101000","000000000000110100","000000000000000000","000000000000001001","000000000000001101","111111111111111001","000000000000011100","000000000000010000","000000000000000001","111111111111110001","000000000000000100","111111111111101011","111111111111101000","111111111111101110","000000000000001111","111111111111101011","000000000000000000","000000000000011001","000000000000000111","000000000000100001","000000000000010010","000000000000000101","000000000000001000","111111111111100000","111111111111110110","111111111111011111","111111111111010011","000000000000000001","000000000000011111","111111111111011110","000000000000100101","111111111110111100","000000000000001111","000000000000001010","111111111111011100","000000000000000101","111111111111110100","000000000000000000","111111111111100011","000000000000000101","000000000000011110","111111111111110010","111111111111001111","111111111111110111","111111111111101010","111111111111110101","000000000000010010","000000000000000011","000000000000001100","000000000000000101","000000000000100010","111111111111111001","000000000000110100","000000000000101010","000000000000000100","000000000000000001","000000000000000111","000000000000000010","000000000000000011","000000000000001100","000000000000000111"),
("000000000000000100","000000000000011100","000000000000010001","000000000000000100","111111111111101101","000000000000000000","000000000000010111","000000000000001101","000000000000001101","000000000000000110","111111111111101011","000000000000111010","111111111111110100","111111111111111010","111111111111110101","111111111111100100","111111111111010111","111111111111100100","111111111111111110","000000000000000010","111111111111110101","111111111111101110","111111111110111111","111111111111011111","111111111111111001","000000000000010010","000000000000000110","000000000000011100","000000000000000111","111111111111100010","000000000000101011","000000000000101101","000000000000001111","000000000000001100","111111111111110100","111111111111111110","000000000000010101","000000000000000011","000000000000001001","000000000000001111","000000000000000000","111111111111100011","111111111111011111","111111111111011001","000000000000001000","000000000000001011","111111111111001101","111111111111110101","000000000000101000","000000000000010001","000000000000000000","000000000000001010","000000000000001100","000000000000001101","000000000000010110","000000000000000101","000000000000101111","000000000000011111","000000000000001001","111111111111110000","000000000000100111","000000000000001100","000000000000010001","111111111111111001","111111111111110111","111111111111110100","111111111111100111","111111111111101001","000000000000101101","000000000000001001","000000000000100000","000000000000000101","111111111111110000","000000000000010101","000000000000000111","000000000000000011","111111111111110110","000000000000010111","000000000000000101","111111111111101001","111111111111011101","000000000000001000","000000000000010001","000000000000000101","000000000000001111","111111111111110000","000000000000001101","000000000000101110","000000000000001000","111111111111111001","111111111111110101","111111111111101100","111111111111011011","111111111111110000","000000000000001101","000000000000000100","111111111111110100","000000000000110011","111111111110010110","111111111111110111","111111111111101111","000000000000001101","000000000000000110","000000000000001000","000000000000001011","000000000000000101","000000000000000111","111111111111111010","111111111111110111","111111111111110100","111111111111111101","111111111111100000","111111111111111111","000000000000100111","000000000000100100","000000000000000101","000000000000100000","000000000000010000","111111111111100111","000000000000010110","000000000000100111","111111111111111111","111111111111110101","111111111111101010","111111111111110101","000000000000010010","000000000000001010","000000000000100100"),
("000000000000011011","000000000000001001","111111111111111111","000000000000010110","111111111111011111","000000000000000011","111111111111111111","000000000000100011","000000000000011001","111111111111111101","000000000000011000","000000000000011001","000000000000100010","111111111111101111","000000000000000011","111111111111101000","111111111111001110","000000000000001110","000000000000000011","111111111111111111","000000000000011000","000000000000000011","111111111111011110","000000000000010101","000000000000010111","000000000000010000","000000000000010101","111111111111111100","111111111111111011","111111111111011011","000000000000110000","000000000000101000","111111111111111101","000000000000000111","000000000000000101","000000000000010100","000000000000000010","000000000000001111","111111111111110001","000000000000000010","111111111111110111","111111111111110010","111111111111110111","111111111111110100","111111111111111000","000000000000000111","111111111110111010","111111111111111000","000000000000001011","000000000000011000","000000000000010011","111111111111100100","000000000000010111","000000000000000100","111111111111111100","000000000000100101","000000000000001100","111111111111110010","111111111111111100","000000000000001010","000000000000011001","000000000000001110","111111111111111101","000000000000000101","000000000000000011","000000000000000110","111111111111010011","111111111111011011","000000000000001100","111111111111111000","111111111111111101","000000000000000111","111111111111110101","000000000000001100","000000000000000001","111111111111111011","000000000000001111","000000000000001110","000000000000011000","111111111111110101","111111111111011001","000000000000011111","000000000000000010","000000000000000000","111111111111111101","111111111111111010","000000000000100111","000000000000100010","111111111111111011","111111111111110010","111111111111111000","111111111111111001","111111111111110110","111111111111101010","000000000000100010","000000000000011000","000000000000010000","000000000000100010","111111111110001110","111111111111101001","111111111111111000","000000000000000111","000000000000001100","000000000000001001","000000000000000111","111111111111111100","000000000000011001","000000000000101010","111111111111110000","000000000000011010","000000000000101001","111111111111100110","000000000000001011","000000000000010000","000000000000101000","000000000000001101","000000000000011100","111111111111101010","000000000000001001","000000000000001000","000000000000011000","111111111111110110","000000000000000100","000000000000100000","111111111111110110","000000000000000101","111111111111111000","000000000000000101"),
("000000000000000000","111111111111101000","000000000000010011","000000000000001001","111111111111101001","111111111111110111","111111111111101101","000000000000111001","000000000000010011","111111111111110111","000000000000000101","000000000000100001","000000000000011010","111111111111011010","000000000000011000","000000000000010101","111111111111011111","000000000000010110","000000000000000101","000000000000001011","000000000000011101","000000000000010100","111111111111110100","111111111111100111","000000000000001011","000000000000000101","000000000000000011","000000000000010101","000000000000000000","111111111111010000","000000000000101010","000000000000001000","000000000000001110","000000000000000000","111111111111110110","111111111111111000","000000000000001011","111111111111110101","000000000000001000","111111111111111001","000000000000000100","111111111111110111","000000000000000010","111111111111110110","111111111111111010","111111111111011101","111111111111010100","000000000000101100","000000000000000011","000000000000000010","000000000000011000","111111111111110110","000000000000001011","000000000000000101","111111111111110110","000000000000000111","000000000000010110","000000000000000010","111111111111111100","111111111111110011","000000000000100000","000000000000000010","000000000000001010","111111111111100111","111111111111101101","000000000000010010","111111111111100110","111111111111110001","000000000000100011","111111111111111001","000000000000001010","000000000000001100","000000000000001110","111111111111100100","111111111111110010","000000000000001000","000000000000010011","111111111111110001","000000000000000100","000000000000001011","111111111111110000","000000000000011001","111111111111111000","000000000000000000","000000000000000000","111111111111110011","000000000000100101","000000000000000010","000000000000000110","111111111111110011","111111111111100100","000000000000001111","111111111111111000","111111111111100011","000000000000000111","000000000000010001","000000000000100001","000000000000111100","111111111110110101","111111111111110000","111111111111111010","000000000000010111","000000000000010001","000000000000000000","111111111111110111","000000000000010000","000000000000001111","000000000000011111","111111111111010011","111111111111111000","000000000000001101","111111111111100001","000000000000001101","000000000000010001","000000000000101110","111111111111100000","000000000000000110","000000000000000101","000000000000000010","000000000000100100","000000000001000000","111111111111100100","111111111111111100","000000000000001100","111111111111111010","000000000000001111","000000000000111000","000000000000000110"),
("000000000000000000","000000000000000101","111111111111110010","000000000000011100","111111111111001110","111111111111111001","111111111111111000","000000000000111001","000000000000010100","111111111111111100","000000000000001000","000000000000100010","000000000000010100","000000000000000111","000000000000010000","000000000000010010","111111111111101110","000000000000000100","000000000000000000","111111111111110110","000000000000010000","000000000000010111","111111111111100001","111111111111001011","000000000000100101","000000000000010111","000000000000001111","000000000000001111","111111111111010010","111111111111000010","000000000000011101","000000000000011011","000000000000100011","111111111111110001","111111111111101001","111111111111101111","000000000000001000","111111111111011111","111111111111110011","111111111111111011","000000000000011100","111111111111000111","111111111111110100","111111111111101100","111111111111111001","111111111111001000","111111111111011011","000000000000001010","000000000000010110","000000000000000101","000000000000011100","111111111111111101","000000000000000010","000000000000000110","111111111111110010","000000000000010100","000000000000000110","111111111111111010","111111111111110101","000000000000000010","000000000000101010","000000000000000100","111111111111111001","111111111111100111","111111111111110000","000000000000000101","111111111111010111","000000000000000000","000000000000100001","000000000000010001","111111111111111111","000000000000000001","000000000000110001","111111111111100101","000000000000001101","000000000000010000","000000000000001110","000000000000000111","000000000000001100","111111111111110001","111111111111101110","000000000000000010","000000000000001000","111111111111011101","111111111111110100","111111111111111001","000000000000010101","000000000000001001","111111111111111010","111111111111100100","111111111111010011","111111111111111111","111111111111111011","111111111111000101","111111111111111001","000000000000010011","000000000000010111","000000000001000101","111111111111000111","111111111111101000","111111111111100011","000000000000000111","000000000000010000","111111111111110110","111111111111110111","000000000000001011","000000000000001101","000000000000011101","000000000000001001","000000000000001101","000000000000100000","111111111111010000","111111111111111101","000000000000000101","000000000000011010","111111111111110110","000000000000011110","111111111111111010","000000000000001000","000000000000011110","000000000000111001","111111111111010110","000000000000000010","000000000000010001","111111111111101100","000000000000100010","000000000000010010","111111111111111100"),
("000000000000001000","111111111111110011","000000000000011111","000000000000000111","111111111111101101","111111111111110001","111111111111101111","000000000000011111","000000000000000000","000000000000000001","111111111111110011","000000000000000000","000000000000010111","000000000000001100","111111111111111101","000000000000010101","111111111111111101","000000000000010111","000000000000011111","000000000000010000","000000000000010011","000000000000110001","111111111111110100","111111111111010111","000000000000011101","000000000000001001","111111111111111010","111111111111111111","111111111111101100","111111111111101010","000000000000100100","000000000000000100","000000000000110101","000000000000010001","000000000000000100","000000000000010111","000000000000001100","111111111111110000","000000000000010110","111111111111110101","000000000000100101","111111111111100100","000000000000001110","000000000000000000","000000000000011010","111111111111011100","111111111111100011","000000000000000111","111111111111111101","000000000000010000","111111111111110110","000000000000001011","111111111111111010","000000000000011011","111111111111110010","000000000000010110","000000000000100101","111111111111011110","111111111111100010","111111111111101010","111111111111110100","000000000000100110","111111111111101010","111111111111110010","000000000000100101","000000000000011001","000000000000000000","111111111111111110","000000000000011110","000000000000000011","000000000000001000","000000000000000110","000000000000110000","000000000000000001","000000000000010100","000000000000001001","000000000000011111","000000000000001011","000000000000000111","111111111111011000","111111111111110001","000000000000010010","111111111111100011","111111111111110001","111111111111100100","111111111111110100","000000000000101001","111111111111100010","000000000000010110","111111111111100100","111111111111111000","000000000000001000","000000000000011110","111111111111001111","000000000000010001","000000000000001111","000000000000000000","000000000000111111","111111111111110011","111111111111100110","111111111111100011","000000000000101001","111111111111111000","000000000000001111","111111111111110011","000000000000001001","000000000000000000","000000000000100010","111111111111110001","000000000000000001","111111111111111111","111111111111001110","000000000000000111","000000000000001000","111111111111111010","111111111111101111","000000000000001111","000000000000000100","111111111111111100","000000000000100101","000000000000110100","111111111111100111","111111111111111011","000000000000011001","111111111111100000","000000000000100001","000000000000011001","000000000000000111"),
("000000000000000101","000000000000001100","000000000000010000","000000000000000010","000000000000010111","111111111111100011","111111111111110101","111111111111111011","000000000000001001","111111111111111000","111111111111100011","111111111111110000","000000000000010111","111111111111111011","000000000000011010","111111111111111010","111111111111110110","111111111111110011","000000000000010001","000000000000000001","000000000000011001","000000000000101101","111111111111100110","111111111111011000","000000000000001110","000000000000010111","111111111111111011","000000000000001000","111111111111111110","111111111111110111","000000000000011010","111111111111111001","000000000000001110","000000000000001100","111111111111111000","000000000000010011","000000000000000000","000000000000001010","000000000000011000","111111111111101100","000000000000001101","111111111111111111","111111111111100110","000000000000000110","000000000000001100","111111111111101011","111111111111100110","111111111111110011","111111111111111101","000000000000000010","111111111111110100","000000000000000101","000000000000001001","000000000000100100","000000000000000000","000000000000000010","000000000000011011","111111111111110001","111111111111101110","000000000000001000","111111111111011110","111111111111101110","111111111111001000","111111111111111001","111111111111111111","000000000000010001","111111111111110000","000000000000001100","000000000000100111","111111111111101000","000000000000011000","000000000000000110","000000000000000010","111111111111110010","000000000000001110","000000000000010101","000000000000010101","000000000000001110","111111111111110011","111111111111001110","111111111111110100","000000000000001100","111111111111011011","111111111111100110","111111111111110001","111111111111111000","000000000000100001","111111111111110100","111111111111111011","111111111111111111","111111111111011010","111111111111110000","000000000000000011","111111111111001101","111111111111110010","111111111111111001","000000000000011000","000000000000110100","000000000000000110","111111111111110001","111111111111111011","000000000000001010","111111111111011111","111111111111110010","000000000000010010","111111111111111100","111111111111111000","000000000000001110","111111111111111010","000000000000001101","111111111111111111","111111111111100001","000000000000001100","000000000000000000","111111111111100101","111111111111001110","000000000000011010","000000000000000000","000000000000000010","000000000000010100","000000000000101001","111111111111010110","000000000000001000","000000000000100001","111111111111100101","000000000000000000","000000000000110001","000000000000011101"),
("000000000000001100","000000000000000010","000000000000001110","000000000000000100","111111111111101101","111111111111001111","000000000000001111","000000000000011001","000000000000000000","000000000000010000","000000000000000010","000000000000001111","111111111111110110","000000000000000101","000000000000000100","111111111111100110","111111111111010010","111111111111101100","000000000000001101","111111111111111010","000000000000010000","000000000001000001","111111111111101100","000000000000000000","000000000000100110","000000000000011111","111111111111011000","000000000000001000","111111111111110110","111111111111110011","000000000000101110","000000000000010101","000000000000110110","111111111111110111","111111111111110101","000000000000001011","000000000000010000","111111111111110110","111111111111111111","111111111111111001","000000000000011000","111111111111111101","000000000000000100","111111111111101010","111111111111110111","111111111111110111","111111111111101101","111111111111011011","000000000000001010","000000000000000000","111111111111011110","111111111111100111","000000000000011001","000000000000110101","000000000000001010","111111111111101110","000000000000011000","000000000000001011","111111111111111111","111111111111110000","111111111111111101","111111111111011000","111111111110111011","111111111111101001","111111111111101111","000000000000011000","111111111111111100","000000000000000001","000000000000011101","000000000000001001","000000000000001101","111111111111111111","000000000000101100","000000000000011000","000000000000101001","000000000000000010","000000000000000110","000000000000011010","111111111111011000","111111111110110101","000000000000000000","000000000000010000","111111111111010000","111111111111011001","000000000000000011","111111111111011010","000000000000011010","111111111111111110","111111111111110110","111111111111111110","111111111111100001","111111111111111110","000000000000000010","111111111111011011","111111111111110011","111111111111111001","000000000000011110","000000000001000111","000000000000110100","111111111111101110","111111111111110110","000000000000001011","000000000000001011","111111111111110000","000000000000001000","111111111111111111","111111111111110100","000000000000010011","000000000000000010","111111111111101101","000000000000010011","111111111111110100","000000000000000011","000000000000100010","111111111111101111","000000000000010011","000000000000011001","000000000000010111","000000000000001000","000000000000110011","000000000000100101","111111111111101111","111111111111111110","000000000000001100","111111111111000011","000000000000000100","111111111111111000","000000000000011011"),
("000000000000100101","000000000000110000","000000000000011111","000000000000100000","111111111111111011","111111111111101101","000000000000000100","000000000000000111","000000000000010010","000000000000001010","111111111111100101","000000000000001011","000000000000000001","000000000000011010","111111111111101111","111111111111011110","111111111111000000","111111111111011011","000000000000000110","111111111111010000","000000000000001000","000000000000100100","111111111111010110","000000000000010001","000000000000010001","000000000000010000","111111111111110100","000000000000100100","111111111111111000","111111111111110111","000000000000100111","000000000000001110","000000000000111001","111111111111111101","000000000000000001","000000000000000011","000000000000000110","111111111111111101","111111111111100110","111111111111110010","000000000000000011","111111111111111101","111111111111110000","111111111111110010","111111111111111100","111111111111110000","111111111111111000","111111111111110010","000000000000001001","111111111111111001","111111111111010011","111111111111100011","111111111111101101","000000000000100101","111111111111111010","111111111111101101","111111111111110110","111111111111111100","111111111111101110","000000000000010010","000000000000000101","111111111111111001","111111111111010111","111111111111110000","111111111111111100","000000000000001000","111111111111011011","111111111111101110","000000000000001100","000000000000000000","000000000000100001","111111111111111000","000000000000100011","000000000000000100","000000000000100001","000000000000100000","000000000000000000","000000000000101011","111111111111111000","111111111111010100","000000000000000001","000000000000110011","111111111111010010","111111111110111110","000000000000000110","111111111111110001","000000000000101011","111111111111111101","111111111111101110","111111111111111011","111111111111110001","111111111111111110","111111111111110000","111111111111101000","111111111111111111","111111111111110000","111111111111101101","000000000001001001","000000000000011000","111111111111110100","000000000000010101","000000000000010100","000000000000001010","000000000000001010","111111111111110100","111111111111111000","000000000000001110","111111111111110101","111111111111101111","111111111111010010","000000000000000111","000000000000011010","000000000000001011","111111111111110111","111111111111101000","000000000000100100","000000000000010010","000000000000000000","111111111111110011","000000000000001101","000000000000010110","111111111111100110","111111111111111010","111111111111110011","111111111111010010","000000000000011000","111111111111111100","000000000000001111"),
("000000000000010101","000000000000010111","000000000000100100","000000000000010101","111111111111110011","111111111111101000","111111111111111101","000000000000001111","111111111111010100","000000000000011010","111111111111010100","000000000000000101","111111111111111001","000000000000110000","000000000000000001","111111111111101110","111111111111001101","111111111111110101","111111111111111000","111111111111101001","000000000000001011","000000000000001001","111111111111101001","111111111111110100","000000000000101011","000000000000000000","111111111111101011","000000000000011001","111111111111010110","000000000000001111","000000000000001001","000000000000010010","000000000000001101","111111111111110011","000000000000000101","000000000000001011","000000000000100100","111111111111111000","000000000000001111","111111111111110101","000000000000000110","000000000000000110","111111111111011000","000000000000000001","111111111111111100","111111111111110100","111111111111001000","111111111111101111","000000000000001010","111111111111011000","111111111111101100","111111111111100100","000000000000000111","000000000000011010","111111111111110001","000000000000000100","111111111111111101","111111111111110011","111111111111110000","111111111111111100","000000000000001100","111111111111101101","111111111111011110","111111111111100100","111111111111110101","000000000000100001","111111111111100001","111111111111101101","000000000000100000","000000000000001110","111111111111111101","111111111111110000","000000000000101100","111111111111111101","000000000000010111","111111111111110111","000000000000100001","000000000000001000","111111111111101100","111111111111011101","111111111111111000","000000000000001010","111111111111001111","111111111111001010","111111111111100101","111111111111111000","000000000000100001","111111111111110010","111111111111100010","111111111111101101","000000000000011001","111111111111111101","000000000000100000","111111111111011111","000000000000000011","111111111111101010","111111111111110111","000000000000001111","000000000000100111","000000000000000011","000000000000001001","111111111111101011","111111111111100010","111111111111101001","111111111111101010","111111111111101011","000000000000100010","111111111111110110","000000000000001011","111111111111111010","000000000000100010","111111111111111110","111111111111111010","000000000000001000","111111111111000011","111111111111110100","000000000000010000","111111111111111000","111111111111111110","111111111111110100","000000000000011010","111111111111100110","111111111111111110","000000000000011001","111111111111101110","000000000000010001","111111111111111000","000000000000101011"),
("000000000000100010","000000000000001111","000000000001000011","111111111111101011","111111111111101111","000000000000000001","111111111111111011","000000000000000101","111111111111001111","000000000000010110","111111111111101111","000000000000100010","111111111111100101","000000000000101010","111111111111111010","111111111111101011","111111111111101000","111111111111110011","111111111111101100","111111111111100101","000000000000001101","000000000000010100","111111111111000000","000000000000000000","000000000000100010","111111111111110000","111111111111111011","111111111111111011","000000000000001010","111111111111101101","000000000000001010","000000000000000000","111111111111111011","000000000000011110","000000000000001100","111111111111101010","000000000000110001","000000000000000010","000000000000010111","000000000000001101","000000000000001000","000000000000100101","111111111111001111","111111111111001101","000000000000011111","000000000000001110","111111111111100100","000000000000010010","000000000000010001","111111111111101010","000000000000001101","000000000000000001","000000000000010001","000000000000010110","111111111111100101","111111111111011110","000000000000010011","111111111111101111","111111111111100111","000000000000010010","000000000000001111","111111111111101110","111111111111110100","111111111111101110","111111111111111101","000000000000101101","111111111111010011","111111111111101111","000000000000011111","000000000000010010","000000000000000010","111111111111110011","000000000000001011","111111111111101001","000000000000001101","000000000000001101","000000000000011111","000000000000010001","111111111111110001","111111111111011011","000000000000011110","000000000000000111","111111111111010011","111111111111001111","000000000000001101","000000000000000101","000000000000010111","000000000000100101","111111111111011101","000000000000001011","000000000000011101","000000000000000100","000000000000011101","111111111111101010","111111111111101101","111111111111111001","111111111111101110","111111111111111001","000000000000011001","000000000000000111","000000000000000000","000000000000001010","111111111111011111","111111111111100101","111111111111101111","111111111111100111","111111111111100111","111111111111101000","000000000000000110","111111111111100010","000000000000000101","000000000000011011","000000000000001001","000000000000001010","111111111111001110","111111111111101010","000000000000001001","111111111111100110","111111111111111100","000000000000001001","000000000000101010","000000000000001011","111111111111101011","111111111111111111","111111111111110010","000000000000100110","111111111111110110","000000000000010011"),
("000000000000110011","000000000000010011","000000000000100111","000000000000010001","000000000000011011","111111111111111111","111111111111110000","000000000000001110","111111111111001101","111111111111110000","111111111111100001","000000000000011111","111111111111010001","000000000000100000","111111111111101101","000000000000001001","000000000000001100","111111111111110011","111111111111111010","111111111111101000","000000000000010110","111111111111011011","111111111111111101","000000000000100101","000000000000001010","111111111111011110","000000000000001111","111111111111111111","000000000000000011","111111111111110011","000000000000011111","111111111111110000","000000000000000000","000000000000000101","000000000000010101","111111111111101010","000000000000001010","000000000000010111","000000000000100100","000000000000011011","000000000000101110","000000000000001101","111111111111011011","111111111111011000","000000000000011010","111111111111111111","111111111111011010","000000000000000110","000000000000001100","111111111111101101","111111111111110011","000000000000001101","000000000000001010","000000000000000010","111111111111101110","111111111111110110","000000000000010100","111111111111110011","111111111111110101","111111111111111110","111111111111101100","111111111111111001","111111111111011110","111111111111011110","000000000000001101","000000000000100010","111111111111100100","000000000000000111","000000000000011101","111111111111111111","111111111111100010","111111111111110101","111111111111111001","111111111111011000","111111111111100100","000000000000001011","000000000000111100","111111111111111101","111111111111100110","111111111111110010","000000000001000001","000000000000100110","111111111111110101","111111111111110110","111111111111111101","000000000000000001","000000000000011101","000000000000101001","111111111111111101","111111111111100100","000000000000011010","000000000000000000","000000000000001110","111111111111111110","111111111111100110","000000000000000110","111111111111010101","000000000000010001","111111111111110100","000000000000001100","000000000000011010","111111111111111001","111111111111101101","000000000000000001","111111111111100111","111111111111010111","000000000000000010","111111111111110011","111111111111111111","111111111111111100","111111111111011111","000000000000011100","000000000000001010","111111111111110011","111111111111010111","000000000000010001","111111111111110111","111111111111011101","000000000000101110","111111111111111110","111111111111110101","111111111111111110","111111111111111001","111111111111011001","111111111111110100","000000000000000110","111111111111101000","000000000000000001"),
("000000000000011110","000000000000000100","000000000000011100","111111111111111110","000000000000001110","111111111111100101","000000000000000000","000000000000000101","111111111111101010","000000000000011011","000000000000000000","000000000000011101","111111111111101000","000000000000100001","111111111111011001","000000000000000111","111111111111110000","000000000000101100","111111111111111100","000000000000010010","000000000000010101","111111111111101011","000000000000001110","111111111111101110","000000000000010100","111111111111110100","000000000000011100","000000000000001101","111111111111111101","000000000000001100","000000000000001010","111111111111111100","000000000000011110","000000000000010001","111111111111110101","111111111111010101","000000000000010001","000000000000011000","000000000000100000","000000000000011010","000000000000100000","000000000000001010","111111111111111001","111111111111010100","000000000000001000","111111111111111100","111111111111111000","111111111111111010","000000000000000000","000000000000000000","000000000000000101","000000000000000001","000000000000011111","000000000000010011","111111111111110111","111111111111100100","000000000000000010","111111111111110011","000000000000000000","000000000000001111","111111111111110001","111111111111110000","111111111111100001","111111111111011011","000000000000000100","000000000000010111","111111111111110010","000000000000000001","000000000000001010","000000000000001001","000000000000000000","000000000000001101","111111111111101110","111111111111011110","000000000000010100","000000000000100110","000000000000001010","111111111111111101","111111111111011011","111111111111101001","000000000000000000","111111111111111100","111111111111111011","111111111111111101","000000000000001011","111111111111101101","000000000000011011","000000000000011001","000000000000000100","000000000000000110","000000000000010001","000000000000010001","000000000000001001","111111111111101110","111111111111110110","111111111111110100","000000000000010011","000000000000010011","000000000000000001","000000000000000111","000000000000001101","111111111111100101","111111111111101001","111111111111110111","111111111111110001","111111111111010100","111111111111111010","111111111111101111","111111111111101101","111111111111111001","111111111111101100","000000000000000100","111111111111111111","111111111111111001","111111111111010110","000000000000000000","111111111111110100","111111111111111110","000000000000001111","000000000000010001","000000000000011101","000000000000011001","111111111111101101","111111111111111000","111111111111101011","000000000000010100","111111111111111110","111111111111101110"),
("111111111111101101","111111111111101110","111111111111111001","000000000000001111","000000000000000001","000000000000001110","000000000000010100","000000000000000011","111111111111111111","111111111111110111","000000000000001011","111111111111011011","000000000000000000","111111111111110001","000000000000010100","000000000000000110","000000000000001100","111111111111110111","000000000000000001","000000000000000001","111111111111101101","111111111111110001","000000000000000101","000000000000001001","111111111111110011","000000000000001111","111111111111111000","000000000000011101","111111111111111100","111111111111111010","111111111111111011","000000000000000110","000000000000011011","000000000000000000","000000000000001110","000000000000000010","000000000000000001","111111111111101110","111111111111111101","111111111111110100","111111111111101010","111111111111111111","000000000000001000","000000000000001001","000000000000000100","000000000000010010","111111111111110100","000000000000000111","111111111111011100","111111111111111010","111111111111111111","111111111111111000","111111111111101011","000000000000000000","111111111111111100","000000000000100010","000000000000000111","000000000000000000","000000000000001010","111111111111110111","000000000000000100","000000000000000101","000000000000001001","000000000000000000","000000000000001011","000000000000000111","000000000000001010","111111111111101110","000000000000000000","000000000000001011","000000000000001100","000000000000001001","111111111111110000","000000000000001011","000000000000001110","000000000000011110","111111111111111111","000000000000100000","000000000000010000","111111111111110001","111111111111111100","000000000000010001","000000000000000111","000000000000000101","000000000000001000","111111111111111111","000000000000010000","000000000000010110","111111111111110010","000000000000010100","111111111111110011","111111111111110011","111111111111111111","111111111111110011","000000000000000000","000000000000000000","111111111111110111","000000000000001100","000000000000010000","111111111111110100","000000000000001011","000000000000000111","000000000000000001","000000000000000100","000000000000001111","111111111111111000","000000000000000101","000000000000000100","000000000000000011","000000000000000010","111111111111110000","000000000000010110","111111111111111011","111111111111111100","111111111111110100","111111111111101110","000000000000001101","111111111111111110","000000000000001100","000000000000010111","111111111111110110","000000000000001000","000000000000001010","111111111111101111","111111111111111101","111111111111111100","111111111111110001","111111111111110111"),
("111111111111101010","111111111111011110","111111111111100101","000000000000011100","000000000000000000","000000000000000011","000000000000001001","000000000000000000","000000000000011011","111111111111111101","000000000000001100","000000000000000000","111111111111110111","111111111111110001","111111111111110110","111111111111111011","000000000000000011","000000000000010011","000000000000000101","000000000000000111","111111111111101000","000000000000001000","111111111111111010","000000000000001011","000000000000001101","000000000000010111","000000000000010110","111111111111111010","000000000000000010","111111111111101111","000000000000000001","111111111111110000","000000000000001101","111111111111111111","000000000000000010","000000000000000101","000000000000011000","000000000000001011","111111111111111000","111111111111110111","000000000000010100","111111111111110010","000000000000011101","000000000000010011","111111111111100111","111111111111101100","000000000000011010","000000000000001001","111111111111111111","111111111111110100","111111111111110010","111111111111111010","000000000000001110","000000000000000010","000000000000010111","000000000000000000","000000000000001011","111111111111110100","111111111111111101","111111111111110111","111111111111110111","000000000000001111","111111111111111000","111111111111101000","111111111111111000","111111111111110101","000000000000000101","000000000000010011","000000000000001101","111111111111101100","000000000000001010","000000000000011100","000000000000001111","111111111111111100","111111111111100110","000000000000010000","000000000000000110","000000000000001101","111111111111101001","000000000000000001","111111111111110001","000000000000000001","000000000000011010","000000000000000001","111111111111110101","111111111111111110","111111111111110101","000000000000001010","000000000000000111","000000000000001011","000000000000001011","000000000000000000","000000000000001101","000000000000001000","111111111111111000","111111111111111001","000000000000000000","111111111111101110","000000000000001101","111111111111110011","000000000000001110","111111111111101111","111111111111101111","000000000000010110","000000000000011000","000000000000001101","111111111111110100","000000000000000010","111111111111111001","111111111111111110","111111111111110100","111111111111110111","000000000000000000","000000000000000000","000000000000001100","000000000000001011","000000000000000000","111111111111101110","111111111111110000","000000000000010011","000000000000011000","000000000000001001","000000000000011000","000000000000001011","000000000000010010","111111111111110110","000000000000000011","111111111111110111"),
("111111111111110101","000000000000010001","000000000000001101","000000000000001010","000000000000001000","000000000000000001","111111111111110011","111111111111101110","000000000000000011","111111111111101100","111111111111110000","000000000000000010","000000000000000011","000000000000001010","111111111111110010","000000000000000101","111111111111111110","111111111111111001","111111111111110001","111111111111111111","000000000000000111","111111111111111001","000000000000001101","111111111111110100","111111111111110000","111111111111110101","000000000000000000","000000000000000011","111111111111111001","111111111111101111","000000000000001100","111111111111110111","000000000000010011","000000000000010001","111111111111101101","111111111111110010","000000000000000000","111111111111110000","000000000000001011","111111111111101100","000000000000000101","111111111111110001","000000000000000111","000000000000001000","000000000000010010","000000000000001011","000000000000000100","111111111111110000","000000000000010100","000000000000000000","111111111111110001","000000000000000100","000000000000001110","000000000000000100","000000000000000010","111111111111110000","111111111111101111","111111111111101101","111111111111110100","000000000000000100","000000000000010000","000000000000001010","000000000000010000","000000000000010000","111111111111110111","000000000000010000","111111111111111001","111111111111110011","000000000000001000","111111111111111000","000000000000001011","000000000000000111","111111111111101101","111111111111101110","111111111111111111","000000000000001110","111111111111110000","111111111111111110","111111111111111000","000000000000000010","000000000000010001","000000000000010010","111111111111101110","000000000000000100","111111111111111000","000000000000000001","000000000000000000","000000000000000000","111111111111110100","000000000000000110","111111111111111010","111111111111110101","000000000000001011","000000000000001011","000000000000000011","000000000000000000","111111111111111110","000000000000010001","111111111111111011","000000000000000000","000000000000001000","111111111111101101","000000000000001011","000000000000000000","000000000000010011","000000000000000000","111111111111110101","000000000000001111","000000000000001101","000000000000000011","111111111111110010","111111111111110101","111111111111110011","000000000000000000","111111111111101100","000000000000000000","000000000000001111","111111111111101110","000000000000001100","111111111111111101","111111111111110011","111111111111110010","111111111111111000","000000000000001010","000000000000001101","111111111111101111","000000000000010000","111111111111111111"),
("111111111111111000","111111111111110111","000000000000000111","000000000000000011","000000000000010001","111111111111111011","111111111111111100","111111111111111010","000000000000010011","000000000000010011","111111111111110101","000000000000000000","000000000000010001","111111111111110111","111111111111110101","111111111111111111","000000000000001000","111111111111111110","000000000000010001","111111111111111010","000000000000010001","000000000000001101","111111111111111101","000000000000001110","000000000000001010","000000000000001111","111111111111111001","000000000000000110","111111111111101101","111111111111101111","111111111111111111","000000000000000011","111111111111111010","000000000000010010","111111111111110100","111111111111111001","000000000000000001","000000000000000100","111111111111111001","000000000000010011","111111111111101110","000000000000001010","111111111111111001","111111111111110101","111111111111110111","111111111111111100","111111111111110011","000000000000000110","000000000000000100","111111111111110001","111111111111110011","111111111111111001","000000000000001000","000000000000001100","000000000000001111","000000000000001000","111111111111111010","000000000000001000","111111111111111000","111111111111101111","000000000000000100","000000000000001001","000000000000000110","111111111111110100","111111111111111110","111111111111111011","111111111111110100","000000000000001111","111111111111111101","111111111111111010","000000000000000111","000000000000001000","000000000000010100","111111111111101101","111111111111110001","000000000000001100","000000000000001010","000000000000000010","111111111111111100","000000000000010100","111111111111101111","111111111111111100","000000000000010010","111111111111110110","000000000000010010","111111111111111011","111111111111110111","000000000000010010","111111111111101101","111111111111101101","000000000000010100","000000000000000100","000000000000000001","000000000000000001","000000000000001011","111111111111111000","000000000000000001","000000000000001000","111111111111101111","111111111111111000","111111111111101111","111111111111110110","111111111111110001","000000000000001111","000000000000000111","000000000000001010","000000000000010001","111111111111110000","000000000000010001","000000000000001010","111111111111110011","111111111111110001","000000000000000001","111111111111111111","111111111111101101","000000000000000101","000000000000010000","111111111111111001","111111111111110011","000000000000010000","000000000000010010","000000000000000011","000000000000001011","000000000000000111","000000000000001110","111111111111110101","111111111111111111","000000000000001100"),
("111111111111111011","000000000000010000","111111111111110101","111111111111110010","000000000000000101","000000000000000001","000000000000000011","000000000000001111","111111111111110011","000000000000010011","111111111111101110","000000000000001000","111111111111111110","111111111111111100","000000000000001000","111111111111101110","111111111111110101","000000000000010010","111111111111111010","111111111111111001","111111111111110011","000000000000001011","111111111111110100","000000000000010001","111111111111110001","000000000000000110","000000000000001011","111111111111111011","111111111111101111","000000000000000111","111111111111101101","000000000000001000","111111111111101111","111111111111110100","000000000000001111","000000000000001010","111111111111110101","000000000000010000","000000000000010010","000000000000010010","000000000000000000","000000000000001010","000000000000000000","111111111111110100","000000000000000001","000000000000001010","111111111111111001","000000000000000000","111111111111110011","000000000000001000","000000000000001010","111111111111101111","111111111111101101","111111111111111111","000000000000000100","000000000000000110","111111111111101111","000000000000001100","111111111111110111","111111111111111111","000000000000010010","000000000000001111","111111111111110001","111111111111110100","000000000000001011","111111111111111010","000000000000001011","000000000000010011","111111111111110110","111111111111110111","111111111111110001","000000000000000100","111111111111111101","111111111111110011","000000000000001100","111111111111111000","111111111111110001","000000000000001000","000000000000001010","000000000000001101","111111111111110010","000000000000001101","000000000000010010","000000000000001000","111111111111110001","111111111111110100","111111111111110100","000000000000000000","000000000000000010","000000000000010010","111111111111111001","000000000000000101","111111111111111111","111111111111111001","000000000000000110","111111111111111011","000000000000001010","111111111111110110","000000000000001110","000000000000001010","111111111111111110","111111111111111001","111111111111110011","000000000000010001","000000000000001110","000000000000010010","000000000000000100","111111111111101110","000000000000010001","111111111111111011","000000000000000001","111111111111110001","000000000000000110","111111111111110111","000000000000000100","111111111111101110","000000000000001000","111111111111101110","111111111111110111","000000000000010100","111111111111111101","111111111111111011","000000000000000110","000000000000001000","111111111111101101","000000000000000111","111111111111111111","111111111111111101"),
("000000000000001100","111111111111111110","111111111111110101","000000000000010010","111111111111111100","111111111111110111","000000000000001010","111111111111111011","111111111111101111","000000000000000101","111111111111111001","000000000000000010","111111111111110010","111111111111110001","000000000000000000","111111111111111110","000000000000000101","000000000000001101","000000000000001011","000000000000000011","111111111111111111","111111111111111100","111111111111111100","000000000000001000","000000000000001010","000000000000001100","000000000000001011","000000000000001000","000000000000000011","000000000000010100","111111111111111000","111111111111110000","000000000000000000","111111111111111111","000000000000000110","111111111111101111","000000000000001101","000000000000010001","111111111111110001","000000000000000110","111111111111110101","000000000000000111","111111111111111111","000000000000001101","111111111111110100","111111111111110101","111111111111111000","000000000000001000","111111111111110100","111111111111111101","000000000000001101","000000000000010010","000000000000010011","111111111111110100","000000000000000000","111111111111110010","000000000000001001","000000000000000011","000000000000010011","111111111111111010","000000000000000100","111111111111110101","000000000000010010","111111111111101100","000000000000010001","000000000000010010","111111111111110001","111111111111110010","111111111111111010","000000000000000010","111111111111111110","111111111111110001","000000000000001111","000000000000000010","000000000000000100","000000000000001011","000000000000000101","111111111111111001","111111111111110110","111111111111111110","111111111111101110","111111111111110110","111111111111111101","000000000000001001","111111111111111111","000000000000001110","111111111111111110","000000000000010100","000000000000000110","000000000000001011","111111111111110101","111111111111111111","000000000000010011","000000000000001111","111111111111111001","111111111111101111","111111111111110101","000000000000010001","111111111111111110","111111111111110001","111111111111101111","000000000000010010","000000000000000111","000000000000000010","000000000000010100","000000000000000111","000000000000001011","111111111111110010","111111111111110000","000000000000000010","111111111111111100","111111111111111001","111111111111110110","111111111111110010","000000000000000011","000000000000010000","111111111111101101","000000000000000000","000000000000001111","111111111111111010","111111111111111110","111111111111101100","000000000000001011","111111111111111111","111111111111110011","111111111111101111","111111111111110110","000000000000001101"),
("111111111111111010","111111111111110001","000000000000000011","111111111111111100","111111111111111011","111111111111110000","000000000000011000","000000000000000000","111111111111111010","111111111111101111","111111111111110111","111111111111101100","000000000000001110","111111111111110111","000000000000000110","000000000000001110","111111111111111101","111111111111111000","000000000000001110","000000000000001001","000000000000001000","000000000000000000","111111111111101111","000000000000001000","111111111111111000","111111111111101110","000000000000000000","000000000000010111","111111111111101010","111111111111111110","000000000000000110","000000000000011000","111111111111111000","111111111111111010","000000000000000101","000000000000010000","111111111111111110","000000000000000010","111111111111110111","000000000000000110","000000000000000000","111111111111111110","000000000000000111","000000000000010001","000000000000001111","000000000000000010","111111111111100111","000000000000010000","000000000000001110","000000000000001001","111111111111110101","111111111111110111","111111111111101111","000000000000000000","000000000000001100","111111111111110101","000000000000000110","111111111111111111","111111111111110010","111111111111110010","000000000000000010","000000000000001011","111111111111100011","111111111111111101","000000000000010110","111111111111111110","000000000000010001","111111111111111001","000000000000001001","111111111111111000","000000000000001010","111111111111101011","000000000000011100","000000000000000010","000000000000001001","000000000000010110","111111111111111000","111111111111111111","111111111111101111","000000000000000000","000000000000010011","000000000000001110","111111111111111011","000000000000000010","111111111111110100","000000000000000010","111111111111111100","000000000000001110","000000000000000011","000000000000000111","000000000000000110","000000000000011011","000000000000000000","000000000000001000","000000000000000111","111111111111111111","111111111111110101","000000000000010011","000000000000000010","111111111111100110","000000000000000100","000000000000000001","111111111111111011","111111111111101100","111111111111111100","111111111111101101","000000000000001010","000000000000000011","000000000000001100","000000000000000000","111111111111110110","000000000000000001","111111111111110111","111111111111111010","111111111111111001","000000000000001001","111111111111110010","000000000000000111","000000000000000111","000000000000000100","111111111111111011","000000000000010001","000000000000001000","000000000000010010","111111111111111001","000000000000010110","000000000000000011","111111111111110010"),
("000000000000011010","000000000000010011","000000000000010100","111111111111110111","000000000000001011","000000000000101111","000000000000010100","000000000000000110","111111111111110100","111111111111101001","111111111111111010","111111111111111101","111111111111010011","111111111111111001","111111111111111100","111111111111100001","111111111111111111","111111111111010110","111111111111100001","111111111111111101","111111111111010101","000000000000000000","000000000000001100","000000000000011000","111111111111110011","000000000000101110","111111111111110100","111111111111111000","000000000000000101","111111111111111111","000000000000011111","000000000000000000","111111111111111111","000000000000000001","111111111111111001","111111111111111110","111111111111101000","111111111111101111","000000000000001010","000000000000000000","000000000000000001","111111111111100000","000000000000001111","000000000000011110","000000000000100000","000000000000000011","111111111111101111","000000000000000101","111111111111011100","111111111111111100","111111111111101010","000000000000011011","111111111111001011","111111111111110011","111111111111100001","000000000000101000","000000000000101001","111111111111011101","111111111111101001","111111111111111100","000000000000001101","111111111111111100","111111111111101111","000000000000011011","000000000000100101","000000000000000110","000000000000001000","000000000000011111","000000000000100001","111111111111101110","000000000000101000","111111111111101001","000000000000001000","111111111111100111","111111111111111010","000000000000010001","000000000000100011","000000000000010010","111111111111101110","111111111111101010","000000000000100100","000000000000110011","000000000000100000","111111111111101010","000000000000010001","000000000000001000","111111111111101111","111111111111110001","000000000000101000","111111111111101111","111111111111110010","000000000000101000","000000000000010111","000000000000010110","000000000000000101","000000000000011011","111111111111111110","000000000000001001","111111111111111011","111111111111100111","000000000000001000","000000000000000010","000000000000011100","111111111111111000","111111111111100010","111111111111111101","000000000000010001","111111111111101011","000000000000100010","111111111111111101","111111111111111111","000000000000010110","000000000000000101","111111111111100111","000000000000001010","000000000000000001","000000000000001011","111111111111101100","000000000000010110","111111111111010111","111111111111111000","000000000000001110","000000000000011101","111111111111010100","111111111111101110","111111111111110010","111111111111100011","000000000000011101"),
("000000000000100110","000000000000001011","000000000000010111","111111111111111100","111111111111111001","000000000000000010","111111111111101010","111111111111110011","111111111111101110","000000000000000010","111111111111110111","000000000000010000","111111111111100010","000000000000001010","111111111111111001","111111111111010010","111111111111110111","111111111111100001","111111111111101111","111111111111110010","111111111111110110","000000000000000001","000000000000010100","000000000000000000","111111111111101101","000000000000001100","111111111111101100","000000000000000000","111111111111011111","111111111111011110","000000000000010010","000000000000000011","000000000000101101","000000000000000010","111111111111101001","111111111111101101","111111111111011100","000000000000000101","000000000000011000","111111111111101110","111111111111010111","111111111111111110","000000000000001011","000000000000000011","000000000000101010","000000000000000000","111111111111101010","111111111111110110","111111111111101110","111111111111101111","111111111111001101","111111111111111001","111111111111010110","000000000000100011","000000000000001101","000000000000100100","000000000000100110","111111111111111010","000000000000000000","000000000000000001","111111111111111011","111111111111110010","111111111110111110","111111111111101110","111111111111101111","111111111111100100","111111111111110010","000000000000000110","111111111111011101","111111111111001111","000000000000101010","111111111111001011","000000000000000000","111111111111111010","000000000000001001","000000000000001011","000000000000010110","000000000000011000","111111111111110111","111111111111011100","000000000000001010","000000000000111010","000000000000001110","111111111111000110","000000000000000010","000000000000000010","000000000000000101","000000000000000000","000000000000001001","000000000000000000","111111111111110000","000000000000101010","000000000000010001","000000000000100000","111111111111111000","000000000000011000","000000000000001000","000000000000100101","111111111111101111","000000000000000011","000000000000010110","000000000000001001","000000000000100000","111111111111101100","111111111111000001","111111111111111110","000000000000011010","111111111111111001","000000000000100101","111111111111111000","000000000000001010","000000000000010100","111111111111110101","111111111111011100","111111111111111010","000000000000010101","000000000000000011","111111111111010011","000000000000110010","111111111111011001","111111111111101001","000000000000010100","111111111111110101","111111111111101110","000000000000000000","000000000000010001","111111111111010001","000000000000111000"),
("000000000000101111","000000000000001101","000000000000010100","111111111111110011","111111111111110001","111111111111110111","111111111111111101","111111111111111000","111111111111111100","000000000000000000","111111111111110010","000000000000000000","111111111111110101","000000000000011111","111111111111111011","111111111111001011","111111111111011110","111111111110111110","111111111111101101","111111111111100101","000000000000000000","000000000000100100","000000000000001011","111111111111110110","111111111111111001","000000000000000100","111111111111101001","111111111111101001","111111111111110001","111111111111110100","000000000000000110","000000000000100111","000000000000010000","000000000000001110","111111111111100100","111111111111011101","111111111111110000","111111111111101010","000000000000001110","111111111111111110","111111111111110000","000000000000000010","000000000000001100","000000000000001000","000000000000011011","111111111111101101","111111111111001000","111111111111101011","111111111111011101","000000000000011001","111111111110101111","111111111111111111","111111111111010010","000000000000011010","000000000000000010","000000000000001110","000000000000101000","111111111111111001","111111111111110100","000000000000010000","000000000000010010","000000000000001100","111111111111011110","111111111111111001","000000000000010111","111111111111110111","111111111111101110","000000000000001011","111111111111011111","111111111111100001","000000000000010100","111111111111100000","000000000000010010","000000000000001101","000000000000010001","000000000000000111","111111111111111110","000000000000001111","111111111111111000","111111111111110101","000000000000010111","000000000000110001","000000000000001100","111111111111001010","111111111111110001","000000000000010100","111111111111100101","111111111111101000","000000000000000011","000000000000000011","111111111111111000","000000000000001011","000000000000001101","000000000000101111","000000000000000101","000000000000110000","111111111111110110","000000000000011111","111111111111101110","000000000000001111","000000000000010101","111111111111111111","000000000000010011","111111111111101000","111111111111010001","111111111111101100","000000000000011110","111111111111100000","000000000001000001","111111111111111000","000000000000010101","000000000000000001","111111111111111000","111111111111111110","000000000000001101","000000000000100000","111111111111111100","111111111111011001","000000000000101101","111111111111101110","111111111111101010","000000000000000101","000000000000011001","111111111111100111","111111111111101011","111111111111110111","111111111111100010","000000000000011110"),
("000000000000101111","000000000000000001","000000000000001110","000000000000011110","111111111111100101","111111111111100010","000000000000101011","111111111111101111","000000000000010001","000000000000001101","000000000000110101","111111111111110000","000000000000000111","000000000000010110","000000000000001001","111111111111011110","111111111111100011","111111111111100011","000000000000001101","111111111111110010","111111111111111101","000000000001011100","000000000000000111","111111111111101010","111111111111110101","111111111111111010","111111111111001100","000000000000001111","111111111111110000","111111111111011110","111111111111111011","000000000000100011","000000000000100010","111111111111110110","111111111111110110","111111111111111110","111111111111101100","111111111111100001","000000000000000000","111111111111110010","111111111111100100","111111111111110101","000000000000001110","000000000000000111","111111111111110001","111111111111111101","111111111111110010","111111111111011111","000000000000000101","000000000001000111","111111111111000100","111111111111001100","000000000000001110","000000000000100111","000000000000100000","000000000000001110","000000000000000011","000000000000010010","000000000000011110","000000000000010011","000000000000011001","111111111111111110","111111111111101001","111111111111111100","000000000000010100","000000000000001101","111111111111100011","000000000000000100","000000000000011110","111111111111010101","000000000000000101","000000000000001000","000000000000001010","000000000000101001","000000000000001000","000000000000000111","111111111111101011","000000000000000111","000000000000011110","111111111111110101","111111111111100101","000000000000001010","111111111111111110","000000000000000111","111111111111101100","000000000000000101","000000000000000000","111111111111110110","000000000000000110","111111111111110111","111111111111110101","000000000000011110","000000000000001110","000000000000001000","000000000000010010","000000000000011111","000000000000010000","000000000000101000","111111111111111010","000000000000100010","000000000000011010","111111111111101111","000000000000011111","111111111111110111","111111111111110001","111111111111111011","000000000000011110","000000000000100101","000000000000100000","111111111111111011","000000000000011111","111111111111111000","111111111111011110","000000000000001000","000000000000011000","000000000000001010","000000000000011110","111111111111110101","000000000000010000","000000000000010111","000000000000001001","111111111111101011","000000000000001100","000000000000001100","111111111111111000","000000000000010000","111111111111101010","000000000000101010"),
("000000000000100101","111111111111111001","000000000000001000","000000000000000011","111111111111110010","111111111111111011","000000000000100100","111111111111011111","000000000000111011","000000000000000001","000000000000010101","111111111111100000","000000000000010100","000000000000011100","111111111111111011","111111111111101011","111111111111001010","000000000000010000","111111111111111011","000000000000011011","000000000000110000","111111111111111011","000000000000101011","000000000000000100","000000000000011010","000000000000011101","111111111110111000","000000000000000100","111111111111111001","111111111111101011","000000000000000111","000000000000100010","111111111111110101","000000000000001010","111111111111101001","111111111111101010","000000000000001101","111111111111110001","000000000000000000","000000000000001000","000000000000010000","000000000000001110","111111111111111000","000000000000001101","111111111111101011","111111111111111100","111111111111011111","111111111111001110","111111111111110101","000000000000110111","111111111111100110","111111111111001100","000000000000011001","000000000000010000","000000000000010011","000000000000010000","111111111111111110","000000000000011101","000000000000100011","000000000000001100","000000000000110101","000000000000001000","000000000000000110","111111111111111101","000000000000000110","000000000000010010","111111111111101011","000000000000000010","111111111111101000","111111111111111100","000000000000011111","000000000000001011","000000000000000000","000000000000100010","000000000000101000","111111111111110000","111111111111100111","000000000000010111","111111111111111110","111111111111111100","111111111111110011","111111111111111111","111111111111101010","111111111111110101","111111111111100001","000000000000001000","000000000000010010","111111111111001111","000000000000001001","000000000000000111","111111111111100010","000000000000000010","111111111111101011","111111111111101101","000000000000011100","111111111111110101","000000000000000010","000000000000010111","000000000000010101","000000000000110001","000000000000000111","000000000000000010","000000000000010011","000000000000000000","000000000000001000","111111111111100101","000000000000101110","000000000000010000","111111111111110101","000000000000000011","000000000000110000","111111111111100010","111111111111110001","000000000000001011","111111111111111000","000000000000011010","000000000000000010","000000000000001110","111111111111110010","000000000000010011","000000000000101010","111111111111100100","000000000000001110","111111111111111101","111111111111011101","111111111111110101","000000000000011001","000000000000000100"),
("000000000000000011","000000000000010101","000000000000101100","000000000000010010","111111111111001111","111111111111011100","000000000000011001","111111111111100001","000000000000101101","111111111111100101","111111111111100100","111111111111011011","000000000000000110","000000000000011101","000000000000011101","111111111111101111","111111111111011110","111111111111101001","000000000000001001","000000000000010010","000000000000010110","111111111111110001","000000000000000010","111111111111111010","000000000000100011","111111111111101001","111111111111001110","000000000000111011","111111111111011110","111111111111110010","111111111111111110","000000000000111100","111111111111110111","111111111111111111","111111111111101010","111111111111111001","000000000000010000","111111111111010101","000000000000001010","000000000000001100","000000000000010011","111111111111011010","111111111111110001","000000000000001111","111111111111011101","111111111111111111","111111111111110010","111111111111100101","000000000000000100","000000000000110100","111111111111100011","111111111111010010","000000000000011011","000000000000101111","000000000000010001","000000000000011101","000000000000010001","000000000000010100","000000000000011111","111111111111111000","000000000001000100","000000000000001011","000000000000011001","000000000000001101","000000000000010100","000000000000000011","111111111111101101","111111111111110001","000000000000000100","111111111111011111","111111111111111100","000000000000011001","000000000000000110","000000000000110101","000000000000111010","111111111111111100","111111111111011000","000000000000010110","000000000000100011","111111111111111011","111111111111110001","000000000000001011","111111111111011110","000000000000000000","111111111111100000","000000000000010110","000000000000001110","111111111111010010","111111111111101111","000000000000001111","111111111111100011","000000000000010101","111111111111111101","111111111111010101","000000000000010101","000000000000000101","111111111111110011","000000000001001011","000000000000101011","000000000000111010","000000000000000101","111111111111100010","000000000000010001","111111111111101010","111111111111111010","111111111111011000","000000000000100111","000000000000010001","000000000000000111","000000000000000001","000000000000110110","111111111111101100","111111111111010111","111111111111101111","111111111111111010","111111111111110111","111111111111111000","111111111111111110","000000000000000011","000000000000101110","000000000000001010","111111111111010100","000000000000011011","111111111111100101","111111111111100100","000000000000000000","000000000000011110","000000000000101100"),
("000000000000000000","000000000000000000","000000000000000100","000000000000000011","111111111111011010","111111111111011101","000000000000101010","000000000000000000","000000000000010000","000000000000000000","111111111111110101","000000000000000010","111111111111101110","000000000000100101","111111111111111010","111111111111110101","111111111111111011","111111111111111101","111111111111100111","111111111111101111","000000000000100011","111111111111110010","000000000000000111","111111111111110000","111111111111111110","000000000000000100","111111111111010101","000000000000111110","111111111111010111","111111111111111001","000000000000010110","000000000001001111","000000000000001100","000000000000000011","111111111111111000","000000000000001100","000000000000010010","111111111111110010","000000000000010100","000000000000000011","000000000000010101","111111111111100011","111111111111010010","000000000000000100","111111111111101000","111111111111101101","111111111111101100","111111111111010000","111111111111101101","000000000000110001","111111111111110011","111111111111110101","111111111111111101","000000000001001011","000000000000100010","000000000000010100","000000000000100101","000000000000111010","000000000000001000","111111111111110110","000000000000101100","000000000000010100","000000000000001110","111111111111100011","000000000000001100","111111111111111011","000000000000000100","111111111111101101","000000000000000111","111111111111101010","000000000000001010","000000000000000110","000000000000010000","000000000000101010","000000000000101010","000000000000011011","111111111111011100","000000000000011101","111111111111111110","111111111111110111","111111111111110001","000000000000011110","111111111111011001","111111111111101101","000000000000000011","111111111111111000","000000000000010110","111111111111011100","000000000000000010","111111111111111110","111111111111100100","000000000000001111","111111111111010101","111111111111001011","111111111111111101","000000000000001111","111111111111111100","000000000000111110","000000000000010111","000000000000110000","000000000000010001","111111111111000011","000000000000001010","111111111111111110","000000000000000101","111111111111101001","000000000000100000","000000000000000101","000000000000101011","111111111111111100","000000000000100101","111111111111110100","111111111111100001","000000000000010011","000000000000010111","111111111111111111","000000000000011010","000000000000000010","000000000000000110","000000000000111010","000000000000000110","111111111111010100","000000000000010110","111111111111101111","000000000000000100","111111111111111011","000000000000001001","000000000000100011"),
("000000000000100100","111111111111100001","000000000000010111","000000000000010111","111111111111111011","000000000000001100","000000000000000110","111111111111101101","000000000000010011","000000000000011100","111111111111111011","000000000000101010","111111111111111011","000000000000100100","111111111111111011","111111111111011011","111111111111010111","111111111111111100","111111111111110100","111111111111101100","000000000000010101","111111111111110011","111111111111101001","111111111111010101","000000000000011111","000000000000010111","111111111111110011","000000000000101000","111111111111110110","111111111111101001","000000000000011000","000000000000111000","000000000000001111","000000000000011101","111111111111111100","111111111111110100","111111111111111011","111111111111110100","000000000000001000","111111111111110111","000000000000011011","111111111111101011","111111111111011111","111111111111111001","000000000000000001","000000000000000011","111111111111111001","111111111111010000","000000000000001001","000000000000011100","111111111111011111","111111111111110011","000000000000010010","000000000000111100","000000000000100001","111111111111100111","000000000000010000","000000000000101100","000000000000001010","111111111111110101","000000000000110100","000000000000010100","111111111111110100","111111111111110000","111111111111111101","000000000000010100","111111111111110000","000000000000000010","000000000000000010","111111111111101001","000000000000001011","000000000000100001","000000000000100001","000000000000011111","000000000000011111","000000000000010010","111111111111100111","000000000000010001","111111111111101000","111111111111011110","000000000000000011","111111111111111110","111111111111001110","111111111111011010","000000000000000101","111111111111110010","000000000000011011","111111111111010100","000000000000000010","111111111111110000","111111111111001100","000000000000010011","000000000000000011","111111111111011101","111111111111110101","000000000000110010","111111111111101101","000000000000111110","000000000000011001","111111111111111001","000000000000101100","111111111111101101","000000000000010101","000000000000010110","111111111111111010","111111111111101111","000000000000000101","000000000000000010","000000000000011100","111111111111101001","000000000000000000","111111111111100011","111111111111111111","000000000000001011","111111111111111111","000000000000010100","000000000000100011","000000000000000000","000000000000010001","000000000001001000","111111111111111000","111111111111111011","000000000000001100","111111111111101101","111111111111110100","000000000000001001","111111111111110100","000000000000010101"),
("000000000000101000","000000000000010100","000000000000011110","000000000000010111","111111111110000000","000000000000010011","000000000000000111","111111111111110101","000000000000000011","000000000000000011","111111111111011101","000000000000100111","111111111111111101","000000000000100110","000000000000010000","000000000000000010","111111111111011010","111111111111101110","000000000000010000","000000000000000001","000000000000010110","111111111111011100","111111111111111100","111111111111110000","000000000000101001","000000000000001001","111111111111110001","000000000000010111","111111111111101010","111111111111110100","000000000000010001","000000000000001111","000000000000111001","000000000000101001","111111111111101100","111111111111100010","000000000000010111","111111111111011100","000000000000001000","000000000000000010","000000000000011110","111111111111101011","000000000000010110","111111111111100010","111111111111110110","111111111111110110","111111111110111000","111111111111011001","000000000000001110","000000000000010100","111111111111101101","111111111111110111","111111111111111110","000000000001000001","000000000000000111","111111111111101110","000000000000100011","000000000000100111","000000000000000100","111111111111101100","000000000001001000","000000000000110011","111111111111111111","000000000000000110","000000000000001000","000000000000101010","000000000000010110","000000000000011011","000000000000010011","000000000000001101","000000000000011011","111111111111110011","000000000001000110","111111111111111001","000000000000010110","000000000000001010","111111111111110000","000000000000010010","111111111111101111","111111111111110000","111111111111111010","000000000000010000","000000000000000001","111111111111000001","111111111111010100","111111111111100111","000000000000001111","111111111111110100","111111111111110000","111111111111001110","111111111111001011","000000000000001101","111111111111110001","111111111111111011","000000000000011111","000000000000001101","000000000000000000","000000000001000000","111111111111100111","111111111111110000","000000000000110110","111111111111110110","111111111111111111","000000000000000100","111111111111111000","111111111111111110","000000000000011100","000000000000001100","000000000000000000","000000000000001100","000000000000000110","111111111111100000","111111111111111100","000000000000001001","111111111111011010","111111111111111000","000000000000100011","111111111111111010","111111111111111111","000000000001000010","000000000000000110","111111111111101000","111111111111111001","111111111111110111","111111111111011000","000000000000001100","111111111111110111","000000000000011000"),
("000000000000010100","000000000000001101","000000000000010111","000000000000010110","111111111110100001","111111111111101111","000000000000001010","111111111111111000","000000000000011011","000000000000010101","111111111111101011","000000000000001110","000000000000011100","000000000000110110","000000000000000000","111111111111110011","111111111110111011","111111111111011111","000000000000010100","000000000000001111","000000000000011101","111111111111110111","111111111111011110","111111111111100100","000000000000100001","111111111111111101","111111111111001000","000000000000100010","111111111111111011","111111111111101011","000000000000101100","000000000000110110","000000000000010100","000000000000101001","000000000000000101","111111111111110000","000000000000001110","111111111111010011","000000000000001100","000000000000001111","000000000000100001","111111111111010001","111111111111111111","111111111111110111","111111111111110010","111111111111111100","111111111111001001","111111111110110111","000000000000010010","000000000000100101","000000000000010010","111111111111100001","000000000000010100","000000000000101111","000000000000001100","111111111111110000","000000000000101110","000000000000111010","000000000000010000","111111111111101100","000000000001010110","000000000001000011","111111111111100010","000000000000001001","111111111111111000","000000000000001101","000000000000000111","000000000000000000","000000000000010111","111111111111110010","111111111111111111","000000000000011001","000000000000111111","000000000000100000","111111111111111111","000000000000010101","111111111111101011","000000000000000011","000000000000011010","111111111111010110","111111111111110110","111111111111111111","111111111111011010","111111111111100011","111111111111110100","000000000000000000","000000000000011011","111111111111011001","000000000000011010","111111111111101111","111111111111010101","111111111111111000","000000000000000000","111111111111100110","000000000000001110","000000000000011100","111111111111111011","000000000001010000","111111111111011110","000000000000000001","000000000000100010","111111111111011101","000000000000011000","111111111111100110","111111111111110011","111111111111101010","000000000000000111","000000000000011101","111111111111111110","000000000000001011","000000000000001111","111111111111110001","111111111111101101","000000000000010100","000000000000010001","000000000000001011","000000000000001000","000000000000000110","111111111111101010","000000000000110110","000000000000000101","111111111111111001","111111111111111011","000000000000000011","111111111111011011","000000000000100101","000000000000001100","000000000000010001"),
("000000000000011010","111111111111011010","000000000000111001","000000000000000101","111111111110110000","111111111111101000","000000000000101000","000000000000000000","000000000000010001","111111111111101111","000000000000000000","111111111111011110","000000000000110000","000000000000110001","000000000000001111","111111111111100111","111111111111001000","111111111111100111","111111111111110101","000000000000010011","000000000000101100","000000000000100011","000000000000000000","111111111111001100","000000000000001111","000000000000010111","111111111110101100","000000000000110011","111111111111011101","111111111111011110","000000000000101010","000000000001011001","000000000000001100","000000000000010011","111111111111101011","000000000000000001","000000000000010011","111111111110110010","000000000000000011","111111111111111000","000000000000011101","111111111111000010","000000000000010101","000000000000001001","111111111111111111","111111111111101111","111111111110101100","111111111111001111","000000000000000100","000000000001000111","111111111111100001","111111111111101000","000000000000000100","000000000001000011","000000000000011111","000000000000011000","000000000000010100","000000000000110111","000000000000100110","111111111111111010","000000000001101000","000000000001001000","000000000000000100","000000000000010000","000000000000011001","000000000000011101","000000000000000110","000000000000010110","000000000000000101","111111111111101011","000000000000000010","111111111111110011","000000000000110100","000000000000101001","000000000000101100","000000000000100101","111111111111110010","000000000000000001","000000000000010001","111111111111110001","111111111111100000","111111111111111110","111111111111110011","111111111111111100","111111111111100011","000000000000000011","000000000000010001","111111111111101100","000000000000000110","111111111111101001","111111111110111000","000000000000100110","000000000000010010","111111111111101010","000000000000101110","000000000000101101","000000000000010010","000000000001000011","111111111111010101","111111111111111000","000000000000001011","111111111111011011","000000000000001101","111111111111110000","111111111111011111","111111111111010111","000000000000110110","000000000000100110","000000000000010100","000000000000011001","000000000000101010","111111111111110110","111111111111001010","111111111111110110","111111111111111101","000000000000001110","000000000000001001","000000000000010111","111111111111110001","000000000000101101","000000000000100101","111111111111010001","000000000000101010","000000000000000000","111111111111011101","000000000000110101","000000000000010001","000000000000101001"),
("000000000000101011","111111111111100101","000000000000101000","111111111111111111","111111111110110100","111111111111101101","000000000000000000","111111111111100001","111111111111110110","000000000000000110","111111111111010100","000000000000001011","000000000000000011","000000000000101000","000000000000011001","111111111111111001","111111111111100100","000000000000000001","111111111111111111","000000000000011001","000000000000111101","000000000000011101","111111111111110010","111111111111110001","000000000000001100","000000000000001111","111111111111100001","000000000000000000","111111111111101010","111111111111011100","000000000000010011","000000000001010001","000000000000011101","111111111111110001","111111111111011110","111111111111100111","000000000000000110","111111111111011000","000000000000010011","000000000000011100","000000000001000000","111111111111100100","111111111111111010","111111111111110000","111111111111110110","111111111111110000","111111111111001101","111111111111101010","000000000000000000","000000000000000111","111111111111111100","111111111111100110","000000000000010101","000000000000111010","000000000000101011","000000000000000101","000000000000000100","000000000000011100","000000000000010010","000000000000000010","000000000001001100","000000000000000111","000000000000000000","111111111111101011","000000000000001011","000000000000000010","000000000000000000","000000000000000111","000000000000110101","000000000000010010","000000000000010100","000000000000010000","000000000001000001","000000000000011010","000000000000110001","000000000000100100","111111111111111110","000000000000011000","000000000000001101","111111111111100110","111111111111111000","111111111111110101","111111111111101111","111111111111111110","111111111111101011","000000000000000001","000000000000011011","111111111111101000","111111111111100111","111111111111111101","111111111111100010","111111111111111101","000000000000001100","111111111111001110","000000000000010010","000000000000000000","000000000000000110","000000000000001111","111111111111101001","111111111111111001","000000000000000110","111111111111110000","000000000000010110","111111111111101010","111111111111011110","111111111110111011","000000000000010011","111111111111111010","111111111111111000","111111111111111111","000000000000011100","111111111111010111","111111111111101000","111111111111110100","111111111111100101","000000000000011110","000000000000000111","000000000000100000","000000000000001110","000000000000111011","000000000000101011","111111111111111101","000000000000001010","000000000000010101","111111111111011100","000000000000011101","000000000000011011","000000000000010000"),
("000000000000111011","000000000000001001","000000000000101001","000000000000000110","111111111110101001","111111111111101011","111111111111111011","111111111111101011","111111111111101011","000000000000010111","111111111111001110","000000000000000111","000000000000001111","000000000001000000","000000000000010001","111111111111111001","111111111111100100","111111111111110010","111111111111100110","000000000000100111","000000000000101101","000000000000001010","111111111111110101","111111111111101011","000000000000011010","000000000000001101","111111111111001001","000000000000010010","111111111111011001","000000000000001001","000000000000011001","000000000001010011","000000000000011111","111111111111101111","111111111111110011","111111111111111110","000000000000010101","111111111111100001","111111111111111101","111111111111111011","000000000000011111","111111111111011111","000000000000000000","111111111111111110","000000000000001100","111111111111111111","111111111111000001","111111111110110100","111111111111110010","000000000000011110","000000000000011011","111111111111011000","000000000000010100","000000000000100010","000000000000010100","111111111111110000","000000000000100111","000000000000011000","111111111111110100","111111111111110010","000000000000101010","000000000000011000","111111111111101101","111111111111101001","000000000000011001","000000000000001111","000000000000010011","000000000000000111","000000000000100100","000000000000000000","000000000000010000","000000000000000001","000000000001010101","000000000000011111","000000000000011001","000000000000011001","111111111111100111","000000000000100101","111111111111101100","111111111111011000","000000000000000001","000000000000001001","111111111111101000","111111111111011101","111111111111011101","111111111111110111","000000000000011100","000000000000000100","000000000000010100","111111111111111100","111111111111010100","000000000000001001","000000000000000100","111111111111101001","000000000000001101","111111111111111101","000000000000001110","000000000000100011","111111111111110000","000000000000100111","000000000000001010","111111111111110000","111111111111111001","000000000000001000","000000000000000000","111111111111010010","000000000000000010","000000000000010011","000000000000011101","000000000000000011","000000000000011111","111111111111001101","111111111111110000","000000000000000111","111111111111101101","111111111111110110","000000000000001001","000000000000011000","000000000000010101","000000000001000011","000000000000001110","111111111111101110","111111111111110111","111111111111110110","111111111111100100","000000000000010010","000000000000100010","000000000000010100"),
("000000000000110100","111111111111111000","000000000000010101","000000000000001111","111111111111011000","111111111111101111","000000000000010111","111111111111011101","000000000000001110","111111111111110100","111111111111011100","000000000000000111","111111111111111100","000000000000101110","000000000000001011","111111111111100100","111111111111101010","111111111111110111","000000000000001100","000000000000010000","000000000000011000","000000000000011011","111111111111101101","111111111111011110","000000000000101001","000000000000000100","111111111111010011","000000000000011000","111111111111100001","111111111111111110","000000000000010010","000000000001100000","000000000000011010","000000000000001101","111111111111110000","000000000000001011","000000000000001010","111111111111111011","000000000000100101","000000000000000001","000000000000101011","111111111111111011","111111111111111011","000000000000011000","111111111111110111","111111111111111111","111111111111011101","111111111111010010","000000000000010000","000000000001000001","111111111111101001","111111111111011101","000000000000000111","000000000001010011","000000000000010110","111111111111110110","000000000000110111","000000000000010111","000000000000001000","111111111111111101","000000000000101101","000000000000100100","111111111111100110","000000000000000000","000000000000101111","111111111111110101","000000000000001010","000000000000111001","000000000000001101","111111111111111011","000000000000001101","000000000000011100","000000000000011110","000000000000011010","000000000000100011","000000000000111100","111111111111100011","000000000000010100","111111111111101101","111111111111010110","000000000000011001","000000000000000010","111111111110111000","111111111111010000","000000000000000010","111111111111110101","000000000000000011","111111111111111010","000000000000101001","000000000000000110","111111111111011010","000000000000011000","000000000000011101","111111111111100000","000000000000001100","000000000000001010","000000000000100000","000000000000101011","111111111111100000","000000000000010001","000000000000001000","111111111111101111","000000000000000001","000000000000001100","111111111111111110","111111111111101111","000000000000100110","000000000000011010","000000000000101111","111111111111100000","000000000000100101","111111111111010100","000000000000000010","000000000000001101","111111111111011111","111111111111111111","000000000000110000","111111111111110100","000000000000100000","000000000000110110","000000000000001001","111111111111110011","111111111111101111","111111111111111000","111111111111001100","000000000000010100","111111111111111101","000000000000101100"),
("000000000000010000","000000000000000100","000000000000010110","000000000000011001","111111111111001011","111111111111100010","000000000000011110","111111111111001101","000000000000011111","000000000000000110","111111111111011011","111111111111100100","000000000000011010","000000000000010010","000000000000010001","111111111111001010","111111111111000011","111111111111110000","000000000000001010","111111111111110111","000000000000101110","000000000000100101","111111111111101111","111111111111100000","000000000000000111","000000000000001101","111111111111001100","000000000000100001","111111111111011110","111111111111101001","000000000000011010","000000000000111011","000000000000010100","000000000000010000","111111111111110000","111111111111110100","000000000000010011","111111111111101001","000000000000010111","111111111111110000","000000000000010001","111111111111100011","000000000000000111","000000000000001001","000000000000000000","111111111111101111","111111111111001000","111111111111010110","000000000000010100","000000000001000010","000000000000001011","111111111111100011","000000000000011011","000000000000101100","000000000000110101","111111111111110111","000000000000001111","000000000000001001","000000000000001010","111111111111110000","000000000000101010","111111111111101000","111111111111101110","000000000000010100","000000000000000010","000000000000000001","000000000000000000","000000000000011110","000000000000001011","111111111111111000","000000000000011011","000000000000011101","000000000000001011","000000000000011100","000000000000001110","000000000000011011","111111111111110111","000000000000000001","000000000000001100","111111111111100110","111111111111111101","111111111111110100","111111111111101010","111111111111011011","111111111111101010","111111111111011100","000000000000000110","111111111111110010","000000000000010010","000000000000011001","111111111111011010","111111111111111011","000000000000000101","111111111111010100","000000000000000000","000000000000001100","000000000000001100","000000000000100001","000000000000010000","000000000000001011","111111111111111011","111111111111110110","000000000000000110","111111111111110101","111111111111100101","111111111111100011","000000000000001111","000000000000100011","000000000000000000","111111111111100110","000000000000101111","111111111111100011","111111111111111011","000000000000001001","111111111111100001","111111111111101001","000000000000101000","000000000000010100","000000000000011001","000000000000101011","000000000000000110","111111111111101110","000000000000010001","000000000000010011","111111111110111100","000000000000011111","000000000000010010","000000000000011000"),
("000000000000010000","111111111111111100","000000000000001110","000000000000010111","111111111111000010","111111111111011001","000000000000000010","111111111111011001","000000000000011010","000000000000100100","111111111111100001","111111111111110110","000000000000011100","000000000000101111","111111111111111110","111111111111100111","111111111111011011","111111111111101010","000000000000100000","000000000000000010","000000000000010111","000000000000111100","111111111111111111","111111111111111110","000000000000001011","111111111111101111","111111111111001010","000000000000001000","111111111111110011","111111111111110110","111111111111111101","000000000000111011","000000000000011011","000000000000010010","111111111111100101","111111111111010010","000000000000010110","111111111111100100","111111111111011111","000000000000010110","000000000001000001","111111111111011001","000000000000010111","000000000000001000","111111111111100011","000000000000001010","111111111111101101","111111111111001110","000000000000000110","000000000000101000","000000000000010011","111111111111100011","000000000000010010","000000000000100011","000000000000100100","111111111111011111","111111111111111000","000000000000101010","000000000000010110","000000000000000011","000000000000001001","111111111111111101","111111111111101011","111111111111101010","000000000000010000","111111111111111001","000000000000011101","111111111111100101","000000000000101001","000000000000100111","111111111111110001","000000000000011111","000000000000001100","000000000000001000","000000000000001000","000000000000001010","111111111111101101","000000000000011101","111111111111111010","111111111111011100","111111111111110100","111111111111101101","111111111111001001","111111111111001001","111111111111100001","000000000000000101","000000000000100101","111111111111111001","000000000000000011","111111111111111100","111111111111011110","111111111111111001","000000000000011101","000000000000010010","000000000000000000","000000000000001101","111111111111100001","000000000000100010","000000000000001000","000000000000101000","000000000000001101","111111111111101000","000000000000000010","111111111111101011","000000000000000011","111111111111011110","111111111111111101","000000000000011111","000000000000000110","111111111111111001","000000000000000010","000000000000000110","111111111111001110","000000000000000110","111111111111011110","111111111111110110","000000000000101111","000000000000111011","111111111111110110","000000000000100100","000000000000011110","111111111111101011","000000000000001100","000000000000011100","111111111111010011","000000000000010111","000000000000001011","111111111111110000"),
("000000000000011100","000000000000010001","000000000000100110","000000000000000110","111111111110110111","111111111111011001","000000000000100000","111111111111111111","000000000000001111","000000000000001001","111111111111001100","111111111111111110","000000000000100111","000000000001010001","000000000000000000","111111111111010111","111111111111000101","111111111111101110","000000000000010111","111111111111101110","000000000000100010","000000000000001011","111111111111001111","111111111111111001","000000000000011001","000000000000010001","111111111111101001","000000000000101000","111111111111101010","111111111111110111","000000000000100010","000000000000101110","000000000000011110","000000000000000010","111111111111100000","111111111111100010","000000000000011101","111111111111011001","000000000000000111","000000000000001011","000000000000100100","111111111111001001","000000000000011000","000000000000000000","111111111111100011","111111111111111110","111111111111100111","111111111111100110","111111111111110000","000000000000100001","111111111111100001","111111111111011000","000000000000001100","000000000000111100","000000000000001011","000000000000001111","000000000000001101","000000000000011100","000000000000010110","000000000000001011","000000000000011011","111111111111111011","111111111111111111","111111111111100111","111111111111110100","000000000000010111","000000000000010101","000000000000000100","000000000000010100","000000000000010001","000000000000001100","000000000000001001","000000000000000000","111111111111111101","000000000000101100","000000000000100111","000000000000000111","000000000000011001","000000000000000001","111111111111011000","111111111111101011","000000000000001100","111111111111011101","111111111111001111","111111111111110110","111111111111011100","000000000000100001","111111111111110111","111111111111110010","000000000000000101","111111111111011100","111111111111111101","000000000000011100","000000000000000100","000000000000011001","111111111111110011","000000000000000000","000000000001000001","111111111111111000","000000000000001101","000000000000010010","111111111111111101","000000000000000100","111111111111110010","111111111111100110","111111111111000110","000000000000100001","000000000000011010","000000000000001111","111111111111010100","000000000000100111","111111111111111111","111111111111110111","111111111111101111","111111111111100011","000000000000010011","000000000000011010","111111111111111000","111111111111110110","000000000000111001","000000000000100000","111111111111100101","111111111111111111","111111111111110101","111111111111011010","000000000000101011","000000000000000111","000000000000011010"),
("000000000000001011","000000000000001001","000000000000101010","000000000000001100","111111111110111011","111111111111101100","000000000000010000","000000000000010011","000000000000000100","000000000000011010","111111111110111010","111111111111011100","000000000000000111","000000000001010010","000000000000100011","111111111111001111","111111111111001010","111111111111111010","111111111111111101","111111111111100011","000000000000110001","000000000000001100","111111111111001100","111111111111111001","000000000000000100","000000000000000010","111111111111011111","000000000000101001","111111111111011001","111111111111110001","000000000000011001","000000000001000110","000000000000001001","111111111111101001","111111111111110001","000000000000010010","111111111111111100","111111111111001100","000000000000001110","000000000000000011","000000000000000111","000000000000000001","000000000000011100","000000000000101000","111111111111101000","000000000000000011","111111111111001011","111111111111101001","111111111111110110","111111111111110001","111111111111110110","111111111111011100","000000000000001001","000000000000101110","000000000000011001","000000000000110001","000000000000001010","111111111111111110","000000000000101110","000000000000000000","000000000000010011","111111111111110000","111111111111101101","000000000000010000","111111111111011110","000000000000111011","000000000000001100","111111111111011000","000000000000010010","000000000000000000","000000000000001100","111111111111100010","111111111111111110","000000000000100010","000000000000110011","000000000000010101","111111111111110011","000000000000100100","000000000000100001","111111111111100010","111111111111110100","000000000000001111","111111111111100001","111111111111001010","111111111111011101","111111111111110110","111111111111111011","000000000000001011","000000000000000100","000000000000000100","111111111111110000","000000000000000000","000000000000000001","111111111111011000","000000000000100111","000000000000001011","000000000000000101","000000000000100011","111111111111111111","000000000000100100","111111111111101100","111111111111100001","111111111111110100","111111111111010111","000000000000001000","111111111110111110","000000000000101011","000000000000010011","000000000000000101","000000000000010110","000000000000011011","111111111111111110","111111111111101110","111111111111110111","000000000000000111","111111111111111010","000000000000010000","000000000000000100","111111111111110101","000000000000011001","000000000000010010","111111111111111001","111111111111111100","111111111111110000","111111111111100011","000000000000010100","000000000000010001","000000000000100111"),
("111111111111110111","111111111111101100","000000000000011011","000000000000001110","111111111111000110","111111111111010101","000000000000011100","000000000000000101","000000000000000011","000000000000011001","111111111111100000","111111111111101010","000000000000011000","000000000000101000","000000000000101000","111111111111111010","111111111111101000","111111111111111001","111111111111111001","111111111111100101","000000000000100100","000000000000101000","111111111111100111","111111111111111001","000000000000010011","111111111111100110","111111111111001101","000000000000100110","111111111111100101","111111111111111011","000000000000001010","000000000000110011","000000000000001011","000000000000000001","000000000000000101","111111111111111010","000000000000000111","111111111111001011","000000000000000001","000000000000000111","000000000000101001","000000000000010101","000000000000001000","111111111111111110","111111111111011011","000000000000001100","111111111111010000","111111111111111110","000000000000001111","000000000000001011","000000000000101110","111111111111101010","000000000000100110","000000000000011011","000000000000010011","000000000000000000","000000000000001001","000000000000000101","000000000000010111","111111111111110000","000000000000101110","111111111111111001","111111111111110110","111111111111111010","000000000000000010","000000000000100011","111111111111110111","000000000000001000","111111111111110010","000000000000111001","000000000000001010","111111111111101101","111111111111010011","000000000000010010","000000000000000101","000000000000001101","111111111111010110","000000000000010001","000000000000000110","111111111111111001","111111111111110111","111111111111101001","111111111111010001","111111111111110100","111111111111100101","111111111111110110","000000000000010000","000000000000000101","111111111111111011","111111111111111000","000000000000001100","111111111111111011","000000000000010100","111111111111110111","000000000000101111","000000000000011000","111111111111111100","000000000000100100","111111111111101101","000000000000110000","111111111111111011","111111111111110001","000000000000000010","111111111111101000","111111111111111011","111111111111011000","000000000000010001","000000000000000111","111111111111111010","000000000000001110","000000000000001110","111111111111111011","111111111111010000","000000000000001111","111111111111111010","111111111111101111","000000000000011111","000000000000010101","111111111111111100","000000000000011000","111111111111110111","000000000000000000","111111111111111111","000000000000010010","000000000000000101","000000000000010011","000000000000000001","000000000000000110"),
("000000000000011011","000000000000011000","111111111111111100","111111111111111010","111111111111000010","111111111111101101","000000000000010101","111111111111101000","111111111111111001","000000000000010010","000000000000000001","111111111111011111","111111111111111110","000000000000100000","000000000000011011","111111111111110010","111111111111111101","000000000000000001","111111111111101011","111111111111110110","000000000000000000","000000000000001011","000000000000010011","000000000000000010","111111111111110110","111111111111111100","111111111111011110","000000000000000010","000000000000001001","111111111111111111","111111111111101110","000000000000010001","000000000000011011","000000000000011111","111111111111100111","111111111111101100","111111111111111100","111111111111110001","000000000000000011","111111111111111100","000000000000001110","000000000000000100","000000000000101000","000000000000010110","111111111111111101","111111111111101101","111111111111101000","111111111111011111","111111111111111010","000000000000010110","000000000000001000","111111111111100000","000000000000001000","000000000000100101","000000000000000001","000000000000010011","000000000000010100","000000000000010011","000000000000110100","111111111111111001","000000000000001100","111111111111111110","000000000000000001","111111111111111111","111111111111101111","000000000000101011","111111111111100100","000000000000100101","111111111111101101","000000000000000001","111111111111111000","111111111111111000","111111111111001101","000000000000010101","000000000000011100","000000000000000001","111111111111100101","000000000000001010","000000000000001100","111111111111100100","111111111111101111","000000000000000000","000000000000010110","111111111111110110","111111111111100101","111111111111101011","000000000000001001","111111111111101011","000000000000011011","000000000000000010","111111111111110000","000000000000100010","111111111111100010","111111111111101010","000000000000101010","000000000000000001","111111111111100110","000000000000011011","111111111111101011","000000000000011100","000000000000100000","111111111111111100","000000000000000001","111111111111011010","111111111111110101","111111111111001101","000000000000101100","111111111111101101","111111111111111000","111111111111110111","000000000000101100","111111111111111111","111111111111111000","000000000000010011","000000000000001011","111111111111111110","111111111111111110","111111111111110000","000000000000010101","000000000000001100","111111111111111001","111111111111111101","000000000000000010","000000000000011000","111111111111101010","000000000000000101","111111111111111010","000000000000100110"),
("000000000000000101","000000000000001010","111111111111110110","111111111111111100","111111111111111001","000000000000001100","000000000000101001","111111111111110010","000000000000010000","000000000000000010","000000000000010001","111111111111011100","000000000000010010","000000000000100001","000000000000001000","111111111111111000","111111111111010101","111111111111110001","111111111111101011","000000000000001110","000000000000000100","000000000000011000","000000000000010011","000000000000010100","111111111111100100","000000000000100101","111111111111011100","000000000000000000","000000000000011001","000000000000001111","111111111111100111","000000000000000110","111111111111101111","111111111111110100","000000000000001000","000000000000010010","111111111111111001","111111111111110100","111111111111111010","000000000000001101","111111111111110101","000000000000010000","000000000000100101","111111111111110101","111111111111110010","000000000000010011","111111111111101110","111111111111010111","111111111111101110","000000000000011010","111111111111010011","111111111111101011","111111111111100000","000000000000011000","000000000000010000","000000000000000110","111111111111111100","111111111111111010","000000000000101010","000000000000001001","000000000000000000","111111111111110101","000000000000001101","000000000000010010","111111111111111000","000000000000011101","111111111111111110","000000000000010001","111111111111011111","111111111111101011","000000000000101100","000000000000000000","000000000000000101","000000000000001111","000000000000011011","000000000000101001","111111111111100000","111111111111110110","000000000000010111","111111111111110000","000000000000000000","000000000000010010","000000000000010010","111111111111101100","111111111111101111","000000000000100101","111111111111110001","111111111111101100","000000000000000111","111111111111101100","111111111111101101","000000000000011111","111111111111011100","000000000000000011","000000000000011001","111111111111110010","000000000000001000","000000000000000111","000000000000000001","111111111111110000","000000000000000011","111111111111110010","111111111111101100","111111111111100101","111111111111111110","111111111111011100","000000000000100010","000000000000010011","000000000000000101","000000000000001011","000000000000010111","000000000000000000","111111111111110001","111111111111110101","000000000000000011","111111111111111011","000000000000010100","111111111111111111","111111111111110011","000000000000001110","000000000000001010","111111111111111100","000000000000001101","111111111111101010","111111111111111010","000000000000001000","000000000000000110","000000000000001000"),
("000000000000001100","111111111111111011","111111111111110111","111111111111110110","111111111111111111","111111111111111101","111111111111111010","000000000000010000","111111111111110111","000000000000000011","111111111111110111","000000000000001111","000000000000000001","000000000000000000","000000000000000000","000000000000010101","111111111111101110","000000000000010000","111111111111111101","000000000000010010","000000000000001001","000000000000000101","000000000000001010","000000000000001110","111111111111111100","111111111111110010","000000000000001001","111111111111110011","111111111111110101","111111111111111000","000000000000000000","000000000000000100","000000000000010000","000000000000000101","000000000000010000","000000000000000000","000000000000001110","111111111111110100","111111111111110101","000000000000000000","000000000000001001","000000000000000000","000000000000001001","111111111111111101","111111111111111001","111111111111110010","111111111111110011","000000000000010000","000000000000000000","111111111111111100","111111111111110111","000000000000000101","000000000000010001","111111111111110101","000000000000001011","000000000000010011","000000000000000000","000000000000000000","111111111111111010","111111111111111010","111111111111111101","000000000000001010","000000000000000101","111111111111111110","111111111111111000","000000000000001011","000000000000001011","111111111111110101","111111111111111110","000000000000011010","111111111111111101","000000000000010010","111111111111101110","000000000000000000","000000000000000100","111111111111111101","111111111111110110","111111111111110111","111111111111110101","000000000000001001","111111111111110110","111111111111110100","000000000000000111","000000000000010111","111111111111111001","000000000000001100","111111111111110110","111111111111111111","000000000000000010","111111111111111010","000000000000000010","000000000000001101","000000000000000001","111111111111101010","000000000000000101","111111111111111011","111111111111111110","111111111111111011","000000000000010100","000000000000010001","000000000000001001","111111111111111000","111111111111101110","000000000000010000","111111111111110100","000000000000010000","000000000000001001","111111111111111000","000000000000001001","000000000000000100","000000000000000111","000000000000000110","111111111111110010","000000000000010100","111111111111110100","111111111111101100","111111111111110100","000000000000001011","000000000000000010","000000000000001111","111111111111110101","000000000000000010","111111111111101101","000000000000001010","000000000000001000","000000000000010001","000000000000010101","111111111111101010"),
("111111111111111100","111111111111110110","000000000000000110","000000000000001011","000000000000000001","000000000000000100","000000000000001111","111111111111110100","000000000000000001","111111111111101111","000000000000000000","111111111111101110","000000000000001011","000000000000000101","111111111111101101","000000000000000000","111111111111110101","111111111111110101","000000000000001010","000000000000000010","000000000000010000","111111111111101110","111111111111110100","000000000000001010","000000000000010011","000000000000000110","111111111111110000","000000000000010001","111111111111111100","000000000000000010","000000000000010000","111111111111111111","111111111111110111","000000000000001111","111111111111110111","111111111111101110","000000000000001100","000000000000010001","000000000000001011","111111111111110011","000000000000001111","111111111111110001","000000000000000110","000000000000000101","111111111111111001","111111111111111011","000000000000000110","111111111111111110","000000000000000111","000000000000001001","111111111111101101","111111111111110001","111111111111101110","000000000000000111","000000000000000110","000000000000000111","000000000000010001","000000000000000001","111111111111111110","111111111111110000","111111111111111010","000000000000000110","000000000000000010","111111111111111001","111111111111111111","000000000000000111","111111111111111011","000000000000000111","000000000000010000","000000000000010001","000000000000001011","000000000000001000","000000000000001110","000000000000001100","111111111111110000","111111111111111000","111111111111111010","000000000000001111","111111111111110111","000000000000010100","000000000000010000","111111111111110111","111111111111101100","111111111111101100","111111111111101111","000000000000001110","000000000000001001","000000000000010010","000000000000000000","000000000000010100","111111111111110100","000000000000010011","111111111111111001","111111111111101110","111111111111101101","111111111111110101","000000000000010010","111111111111101110","111111111111111110","000000000000001110","000000000000000100","000000000000001010","000000000000000000","000000000000001000","111111111111110001","000000000000000101","000000000000000100","111111111111110010","000000000000000110","111111111111110110","000000000000000000","111111111111111101","111111111111110101","000000000000000000","000000000000001001","111111111111110100","000000000000001100","000000000000000100","000000000000001000","111111111111110111","000000000000001001","111111111111110110","111111111111110000","000000000000001100","111111111111101101","111111111111110101","111111111111111100","000000000000010000"),
("000000000000010001","000000000000001010","000000000000000111","111111111111101101","000000000000001100","111111111111111101","000000000000001011","000000000000010011","000000000000001110","111111111111110000","000000000000001100","111111111111110101","111111111111110011","000000000000001100","000000000000001010","111111111111111100","111111111111111010","000000000000010010","111111111111110100","000000000000001100","111111111111110111","111111111111111000","000000000000010011","111111111111110000","000000000000001110","111111111111111011","111111111111110110","000000000000010011","000000000000010100","111111111111111001","111111111111110111","000000000000010000","111111111111110101","111111111111111110","111111111111110111","000000000000010100","000000000000001000","000000000000010000","000000000000010010","000000000000010000","000000000000010000","111111111111110000","111111111111111011","111111111111111100","111111111111101110","111111111111111010","111111111111101110","111111111111111111","000000000000000010","111111111111110011","000000000000001111","000000000000001100","000000000000000011","000000000000010001","111111111111111010","000000000000000011","000000000000001010","000000000000001111","111111111111111101","000000000000000110","111111111111110001","111111111111110010","000000000000001001","111111111111111011","000000000000000111","111111111111101101","000000000000010001","111111111111111001","000000000000001111","000000000000001100","000000000000001100","111111111111111100","000000000000000010","000000000000001011","000000000000010001","000000000000000000","111111111111111111","111111111111101110","000000000000001011","111111111111110010","111111111111110000","111111111111111100","111111111111111101","111111111111111011","111111111111110000","111111111111110100","111111111111110011","000000000000000000","000000000000010011","000000000000001001","000000000000001100","000000000000000101","000000000000001101","000000000000010010","111111111111111111","000000000000010001","000000000000000100","000000000000000000","111111111111110001","000000000000010001","000000000000001100","111111111111110001","000000000000001000","111111111111101111","111111111111110101","111111111111101111","000000000000000000","000000000000001010","111111111111110000","111111111111110000","000000000000001101","000000000000010000","111111111111111011","111111111111111110","000000000000000000","000000000000001010","111111111111110001","000000000000000011","000000000000000010","111111111111101110","000000000000010010","111111111111101110","111111111111110101","111111111111111111","111111111111101101","111111111111111110","000000000000010100","111111111111111001"),
("111111111111110111","111111111111110011","111111111111111101","111111111111111001","111111111111101111","111111111111111111","111111111111110110","111111111111110101","000000000000000111","000000000000001111","111111111111110110","111111111111101111","000000000000000101","000000000000010010","000000000000010010","111111111111111011","111111111111110001","000000000000010001","000000000000000011","111111111111111000","111111111111110100","111111111111101111","111111111111111001","111111111111101100","111111111111110010","000000000000001101","000000000000000010","111111111111110011","111111111111110001","000000000000001011","111111111111110000","000000000000000000","111111111111111011","111111111111111100","000000000000001100","000000000000001100","000000000000010000","111111111111110100","000000000000001100","111111111111110011","000000000000001001","111111111111111000","000000000000000111","111111111111111001","111111111111111010","111111111111101111","000000000000010000","111111111111101111","111111111111101101","111111111111110000","111111111111111010","111111111111101110","111111111111111010","111111111111111010","111111111111111111","111111111111110111","000000000000010000","111111111111111010","111111111111110110","000000000000000000","000000000000000110","000000000000010001","111111111111111111","000000000000000100","111111111111110111","000000000000001100","111111111111111110","000000000000001001","111111111111111101","000000000000010001","111111111111110111","000000000000001010","000000000000001011","000000000000010010","000000000000001001","111111111111111010","111111111111110101","111111111111111110","000000000000010010","111111111111110001","111111111111110101","111111111111111100","000000000000001101","111111111111101101","000000000000000100","000000000000001010","000000000000010001","111111111111110011","000000000000000100","111111111111110001","000000000000001100","111111111111110001","000000000000001001","111111111111110000","111111111111110110","000000000000001011","000000000000010001","000000000000000010","000000000000000101","111111111111101100","000000000000001111","000000000000010010","000000000000000001","111111111111110100","000000000000000110","000000000000010011","111111111111110101","111111111111111011","000000000000000001","111111111111111011","111111111111110000","000000000000001110","000000000000000100","111111111111101100","111111111111110001","000000000000000000","000000000000010001","111111111111110111","000000000000000100","000000000000000101","000000000000010011","000000000000001010","111111111111111101","111111111111111010","111111111111101111","111111111111111110","111111111111101110","000000000000000001"),
("000000000000001010","000000000000000000","000000000000001010","111111111111110110","000000000000000000","000000000000000000","000000000000010010","000000000000001100","111111111111101110","111111111111111011","000000000000010000","000000000000010000","000000000000000101","000000000000001111","000000000000000100","000000000000001110","111111111111101101","111111111111110001","000000000000001101","000000000000001011","000000000000001111","000000000000000011","000000000000001111","111111111111110111","000000000000000000","111111111111111111","111111111111110001","000000000000000101","000000000000010010","000000000000010000","000000000000001000","111111111111110100","000000000000001001","000000000000001110","111111111111111111","000000000000001110","000000000000000010","111111111111110110","000000000000000000","000000000000001001","111111111111111001","111111111111110000","111111111111110111","111111111111110101","000000000000000001","111111111111101101","000000000000000110","111111111111111001","000000000000001111","111111111111111110","111111111111111111","111111111111111011","111111111111111001","000000000000001001","111111111111111110","000000000000001010","000000000000000011","000000000000000110","000000000000001100","111111111111111110","111111111111110100","111111111111111100","000000000000001100","000000000000010011","111111111111101100","000000000000001011","111111111111110011","000000000000000011","111111111111110100","000000000000001000","111111111111111101","000000000000010100","111111111111110100","000000000000000101","000000000000000001","111111111111110111","000000000000000100","000000000000000101","000000000000010010","000000000000000000","111111111111111110","000000000000001000","000000000000001100","000000000000010011","111111111111110011","000000000000001101","111111111111101100","111111111111111000","111111111111111011","000000000000001101","000000000000000110","000000000000010010","111111111111110100","111111111111110101","111111111111110011","111111111111110010","000000000000001010","000000000000000101","000000000000001001","000000000000010100","111111111111101110","000000000000001110","000000000000010000","000000000000001000","000000000000000000","000000000000010000","111111111111111011","000000000000001101","111111111111111000","111111111111111100","000000000000010100","000000000000000000","000000000000000011","000000000000001101","111111111111111001","000000000000000011","111111111111101111","111111111111111110","000000000000000101","111111111111110000","111111111111110111","000000000000001011","111111111111111000","000000000000001101","000000000000000110","111111111111101100","111111111111110111","000000000000010011"),
("111111111111111001","000000000000001010","000000000000001110","000000000000001100","000000000000010001","000000000000000011","000000000000000001","111111111111111010","000000000000010011","111111111111110111","000000000000010011","000000000000001001","000000000000000111","000000000000010011","000000000000010010","000000000000010001","111111111111110100","111111111111111101","111111111111110001","111111111111110010","111111111111110111","000000000000010001","111111111111101100","000000000000000101","000000000000000100","111111111111101100","111111111111101101","000000000000000110","111111111111110000","000000000000010000","000000000000010010","111111111111111111","000000000000000100","000000000000000001","111111111111110111","111111111111111001","111111111111110110","000000000000001000","111111111111110001","111111111111101111","111111111111110100","000000000000000010","000000000000001001","111111111111101101","000000000000000010","000000000000000000","111111111111101110","000000000000001011","111111111111110111","000000000000001111","111111111111101111","000000000000010001","000000000000000001","000000000000001011","111111111111101111","000000000000001010","000000000000001101","000000000000000100","111111111111111110","000000000000000111","111111111111110001","111111111111110100","111111111111110111","000000000000000101","111111111111110011","111111111111111010","000000000000010100","111111111111111011","111111111111101100","111111111111111001","111111111111101100","111111111111110101","111111111111110001","000000000000000000","111111111111110100","000000000000000010","111111111111110010","111111111111111000","111111111111110101","000000000000000001","111111111111101101","000000000000000111","000000000000010001","000000000000001101","000000000000000010","000000000000000000","111111111111111011","111111111111101111","000000000000000000","111111111111111101","000000000000001010","000000000000001101","111111111111110011","000000000000001100","000000000000001001","000000000000000011","000000000000000101","000000000000001011","111111111111101101","111111111111111111","111111111111110000","000000000000001100","111111111111111110","111111111111111111","111111111111111000","000000000000010000","000000000000001011","111111111111110000","000000000000000000","111111111111111011","000000000000001001","000000000000010001","111111111111101100","111111111111101101","000000000000001101","000000000000000010","111111111111111000","111111111111110001","111111111111110011","111111111111101110","111111111111111100","000000000000001101","000000000000001111","000000000000000110","111111111111110010","000000000000000110","111111111111110100","111111111111111110"),
("111111111111111110","111111111111111111","000000000000000001","111111111111110110","000000000000000111","111111111111101111","000000000000000110","000000000000000000","111111111111110010","000000000000000110","000000000000001001","111111111111110011","111111111111111100","000000000000001010","111111111111111100","000000000000001011","000000000000000011","111111111111111000","111111111111110011","111111111111111111","000000000000001110","000000000000000110","111111111111111011","111111111111111111","000000000000000111","111111111111110010","111111111111101100","000000000000001011","000000000000000000","000000000000000101","000000000000000010","000000000000000111","111111111111110011","111111111111110000","111111111111110101","111111111111101111","000000000000000100","000000000000001000","111111111111111110","111111111111111011","111111111111110111","111111111111111100","000000000000000110","000000000000000010","000000000000010000","111111111111111000","111111111111111110","111111111111101111","111111111111110101","000000000000000111","111111111111111010","000000000000000010","111111111111111011","111111111111111100","111111111111111111","111111111111110010","000000000000000101","000000000000001010","111111111111110001","000000000000000000","000000000000001111","111111111111111010","111111111111111110","000000000000001010","111111111111101111","111111111111111011","111111111111110111","000000000000000011","111111111111111100","111111111111110000","000000000000010010","111111111111111100","000000000000001100","000000000000000011","000000000000000101","000000000000000100","000000000000001010","000000000000010001","000000000000010010","000000000000001001","000000000000010001","000000000000010011","111111111111101111","111111111111111010","000000000000010001","111111111111101110","000000000000010100","111111111111111110","111111111111110100","111111111111110010","000000000000010001","111111111111111101","000000000000001011","000000000000001011","111111111111110001","000000000000010100","111111111111110010","111111111111111111","111111111111110101","000000000000001001","111111111111110010","000000000000010011","111111111111110111","000000000000000001","111111111111110101","000000000000010100","000000000000010000","111111111111110110","111111111111101101","000000000000010001","111111111111110101","000000000000001111","111111111111110110","111111111111111001","000000000000010010","111111111111111000","000000000000000011","111111111111110100","111111111111110000","111111111111110101","000000000000001111","111111111111110011","000000000000010000","111111111111110000","000000000000001101","000000000000000111","000000000000001110","111111111111110001"),
("000000000000001101","000000000000001111","111111111111110001","000000000000000101","000000000000000110","111111111111110100","111111111111100011","000000000000001101","111111111111110101","000000000000001010","000000000000010001","111111111111111001","000000000000000000","111111111111100100","111111111111110001","111111111111101110","111111111111111100","000000000000000000","000000000000000110","111111111111110101","000000000000001000","000000000000001100","000000000000000001","111111111111110111","111111111111110110","111111111111111110","000000000000010110","111111111111100001","000000000000000011","111111111111110011","111111111111111010","000000000000001100","111111111111111000","111111111111110011","000000000000100000","000000000000010001","000000000000001011","000000000000011010","000000000000000011","000000000000010111","000000000000001111","111111111111111011","000000000000000010","111111111111111110","111111111111110001","111111111111110000","000000000000000001","111111111111111000","000000000000010011","000000000000010001","000000000000001100","000000000000001011","000000000000011000","111111111111101101","111111111111111111","111111111111111111","000000000000010000","000000000000001000","111111111111111111","000000000000001111","111111111111101000","000000000000001011","111111111111111001","111111111111110110","111111111111110111","000000000000010001","111111111111110101","111111111111110101","000000000000001010","000000000000000001","111111111111111110","000000000000001110","111111111111111101","111111111111111010","111111111111101111","000000000000001000","111111111111101011","111111111111100001","000000000000001000","000000000000001110","000000000000000001","111111111111101010","000000000000000000","000000000000011110","000000000000000001","000000000000001010","111111111111110011","000000000000001100","111111111111111011","111111111111111100","000000000000000000","111111111111111000","000000000000001000","111111111111111000","111111111111100101","000000000000000000","111111111111111110","111111111111100100","111111111111110111","000000000000010000","111111111111110110","000000000000000000","111111111111101010","111111111111101100","000000000000000000","000000000000000110","111111111111100101","000000000000001110","111111111111101110","111111111111110011","111111111111101010","000000000000000101","111111111111110110","000000000000011100","111111111111111000","111111111111100100","111111111111111101","000000000000000110","111111111111101001","000000000000000010","000000000000010110","000000000000001100","111111111111111010","000000000000001001","000000000000011110","111111111111101111","111111111111110111","111111111111100000"),
("111111111111101111","111111111111111001","000000000000000100","111111111111110011","111111111111111011","000000000000000000","111111111111100110","000000000000001100","111111111111110001","000000000000000100","000000000000011100","111111111111110101","111111111111111101","111111111111101011","000000000000010111","111111111111110101","111111111111110100","000000000000010001","000000000000011010","000000000000010011","111111111111111011","000000000000010011","000000000000010001","111111111111110010","000000000000000100","111111111111110000","111111111111111100","111111111111100011","000000000000010100","111111111111110000","111111111111110100","000000000000001110","111111111111111010","000000000000010010","000000000000010101","111111111111110100","000000000000010100","000000000000100000","111111111111111011","000000000000000100","000000000000000000","000000000000000000","000000000000010000","111111111111110111","111111111111101001","111111111111110100","000000000000010011","111111111111101111","000000000000010011","111111111111111011","000000000000000110","111111111111111011","111111111111111101","111111111111111110","111111111111110010","000000000000001101","111111111111110000","111111111111111001","000000000000000000","000000000000000100","111111111111111110","000000000000001000","000000000000010000","000000000000000001","000000000000000111","111111111111110100","111111111111100101","111111111111110011","000000000000001111","000000000000100100","111111111111101100","000000000000000111","111111111111111000","000000000000001000","000000000000001001","111111111111100000","111111111111110010","111111111111111001","000000000000000110","000000000000010010","000000000000001010","111111111111100111","111111111111101110","000000000000010001","000000000000001011","000000000000001100","111111111111111111","111111111111110110","000000000000001011","000000000000001011","111111111111111000","111111111111111101","000000000000001110","000000000000001000","000000000000000000","111111111111101100","111111111111111101","111111111111110101","111111111111110000","000000000000011111","111111111111110000","111111111111101011","000000000000000011","111111111111100000","000000000000001001","111111111111111010","111111111111100010","000000000000010101","111111111111011100","111111111111111100","111111111111101010","111111111111111010","111111111111100010","000000000000010110","000000000000000001","000000000000000001","111111111111100111","000000000000000100","111111111111101100","000000000000000101","111111111111111110","000000000000001011","000000000000001111","000000000000101110","000000000000010111","111111111111110101","111111111111111100","111111111111100101"),
("000000000000000101","111111111111101110","000000000000010010","111111111111011110","111111111111111011","111111111111101111","000000000000000111","111111111111110001","000000000000000000","111111111111111111","000000000000111111","111111111111110100","000000000000011010","000000000000100001","111111111111111000","000000000000010100","111111111111111010","000000000000100100","000000000000010001","111111111111111101","000000000000000101","000000000000100100","000000000000010001","111111111111110101","000000000000000011","000000000000000111","111111111111101010","111111111111111010","111111111111111100","111111111111111001","000000000000000100","000000000000011001","111111111111111100","000000000000001000","000000000000010101","111111111111100110","111111111111111100","111111111111110000","111111111111100111","111111111111110000","000000000000011010","000000000000010001","000000000000011111","000000000000000011","111111111111100000","111111111111101111","000000000000010010","000000000000001001","111111111111111010","000000000000000010","111111111111110000","111111111111110100","000000000000000100","000000000000010000","000000000000000110","000000000000001001","111111111111111111","000000000000101000","000000000000001011","111111111111101101","000000000000001101","000000000000000110","000000000000001101","111111111111101010","111111111111111101","000000000000011100","111111111111111100","000000000000001001","000000000000001101","000000000000000000","000000000000000111","000000000000001110","111111111111110110","000000000000000101","111111111111111110","111111111111110110","111111111111100110","111111111111101111","111111111111111010","111111111111100100","111111111111100110","111111111111110011","111111111111100000","000000000000000000","111111111111101001","111111111111110011","111111111111110100","000000000000001011","111111111111110011","111111111111111101","111111111111111011","000000000000000011","000000000000101000","111111111111111101","000000000000010011","000000000000000101","111111111111111110","000000000000001011","000000000000000111","000000000000011001","000000000000001101","000000000000000100","000000000000011011","111111111111011101","111111111111111000","111111111111110100","000000000000010010","000000000000000110","111111111111101001","000000000000001011","000000000000100010","111111111111101101","111111111111100110","111111111111110011","000000000000000000","000000000000000111","000000000000000011","000000000000011011","111111111111111001","000000000000001111","000000000000000110","111111111111111011","111111111111111100","000000000000100111","111111111111101101","111111111111111100","000000000000000110","000000000000001010"),
("000000000000101000","000000000000000000","000000000000010111","111111111111101001","000000000000000100","111111111111111010","000000000000011101","111111111111101101","000000000000000000","111111111111110011","000000000000111011","000000000000000101","000000000000001000","000000000000101000","000000000000001111","111111111111111010","111111111111100110","000000000000000001","000000000000001110","000000000000000111","000000000000001011","000000000000010010","000000000000110101","111111111111110000","000000000000100001","000000000000001010","111111111111111000","000000000000010010","111111111111110101","000000000000000101","111111111111111100","000000000000011001","000000000000010011","111111111111111110","111111111111101111","000000000000000111","000000000000001110","111111111111111000","111111111111111001","111111111111110001","000000000000001001","111111111111111010","111111111111111110","000000000000000101","111111111111101011","111111111111110011","111111111111110100","111111111111110101","111111111111111111","000000000000011110","111111111111101111","111111111111111101","111111111111110100","111111111111111011","000000000000001111","000000000000000001","000000000000001100","000000000000100110","111111111111111110","000000000000001000","000000000000001101","000000000000010010","000000000000001000","000000000000000111","111111111111011010","000000000000100100","000000000000000111","111111111111111001","000000000000010010","000000000000001100","111111111111111010","000000000000001111","000000000000001101","000000000000001000","111111111111111011","000000000000010010","000000000000000110","000000000000001011","000000000000000010","111111111111111111","000000000000001011","000000000000000011","111111111111101000","000000000000010100","000000000000000010","111111111111111100","111111111111110100","111111111111101100","111111111111110010","111111111111101110","111111111111111001","000000000000000001","000000000000001001","000000000000011010","000000000000011001","111111111111110110","111111111111111110","000000000000001011","000000000000000000","111111111111111001","000000000000011000","111111111111011110","000000000000001100","000000000000001011","111111111111100010","111111111111110000","000000000000000001","000000000000000111","111111111111101000","111111111111110000","000000000000010110","000000000000000000","111111111111101001","000000000000000110","000000000000001101","000000000000010100","111111111111101110","000000000000010110","111111111111110111","000000000000000010","000000000000001111","111111111111110010","000000000000000010","000000000000001000","111111111111111011","111111111111110100","000000000000010000","111111111111111011"),
("000000000000010011","111111111111110110","111111111111111010","111111111111111111","111111111111100011","111111111111110001","000000000000100010","111111111111101100","000000000000000001","111111111111100111","000000000001000100","000000000000000011","111111111111111100","000000000000100001","000000000000010101","000000000000000011","111111111111011001","111111111111110100","000000000000011001","111111111111111010","000000000000011000","000000000000001111","000000000000011000","000000000000000111","000000000000100010","000000000000011000","111111111111100111","000000000000011100","111111111111100110","000000000000010101","111111111111110011","000000000000000011","000000000000001000","000000000000000000","000000000000001110","000000000000000110","000000000000001000","111111111111101000","000000000000000000","111111111111101001","000000000000010101","000000000000001000","111111111111111111","000000000000011011","111111111111100111","000000000000000010","000000000000011100","111111111111011110","111111111111101100","000000000000010100","111111111111011101","111111111111100000","000000000000011001","111111111111110010","000000000000000010","111111111111111001","000000000000010001","000000000000010011","000000000000100010","111111111111110100","000000000000010011","000000000000000100","111111111111111111","000000000000000001","111111111111111010","000000000000010001","000000000000011001","111111111111111001","000000000000001111","000000000000001110","111111111111110001","111111111111111100","000000000000100110","000000000000011000","111111111111101001","000000000000001110","111111111111101011","111111111111110110","111111111111110010","000000000000000100","000000000000000000","111111111111110111","000000000000000001","111111111111111000","111111111111111000","000000000000000100","000000000000000100","111111111111100111","111111111111111110","111111111111110100","111111111111100000","000000000000001101","000000000000001101","000000000000000100","000000000000011010","111111111111110110","000000000000000000","000000000000010010","111111111111111001","111111111111110011","000000000000001001","000000000000000011","000000000000010010","111111111111101110","111111111111101110","111111111111011100","000000000000000010","000000000000010010","111111111111101010","111111111111101100","000000000000010011","111111111111101110","111111111111110111","000000000000001000","111111111111100001","000000000000001111","111111111111111010","000000000000000101","000000000000001011","000000000000000000","111111111111110111","111111111111111110","000000000000000111","000000000000001110","111111111111101101","000000000000000000","000000000000010110","111111111111110110"),
("111111111111111010","111111111111101001","111111111111111000","111111111111111111","111111111111111101","111111111111101001","000000000000011100","000000000000000001","111111111111111010","111111111111111101","000000000000110100","000000000000000011","000000000000010101","000000000000110101","111111111111111000","000000000000010011","111111111111110011","000000000000000000","000000000000000100","111111111111111000","000000000000100111","000000000000010000","000000000000000001","111111111111110110","000000000000001000","111111111111111101","111111111111110101","111111111111111000","000000000000000000","111111111111110011","111111111111110010","000000000000010101","000000000000001100","000000000000001101","000000000000010001","111111111111111101","000000000000001000","111111111111110010","000000000000001001","111111111111111001","000000000000100011","000000000000010000","000000000000000100","000000000000010100","111111111111110110","111111111111111001","000000000000100010","111111111111101111","111111111111110111","000000000000010100","111111111111100010","111111111111110000","000000000000001110","111111111111110110","000000000000000001","000000000000010000","000000000000010000","000000000000000110","000000000000010100","000000000000001011","000000000000000111","000000000000010001","111111111111110111","000000000000001100","111111111111111001","000000000000100000","000000000000000111","111111111111101010","000000000000101101","000000000000010001","000000000000000100","111111111111111100","000000000000001001","000000000000010011","111111111111110000","111111111111111101","111111111111100100","000000000000000100","000000000000010100","000000000000000000","111111111111110100","000000000000001001","000000000000000000","000000000000000011","111111111111101001","000000000000011000","111111111111111110","111111111111100101","111111111111101110","111111111111101110","111111111111110110","111111111111101111","000000000000110100","000000000000001001","000000000000010101","111111111111111011","111111111111111011","111111111111111101","111111111111111111","111111111111111101","000000000000010010","111111111111010100","000000000000001110","111111111111110101","111111111111111000","111111111111011101","111111111111111000","111111111111111110","111111111111101001","000000000000000011","000000000000011110","111111111111110000","111111111111101011","000000000000000000","111111111111111110","000000000000001101","000000000000000110","000000000000000010","111111111111101101","000000000000000011","000000000000000000","111111111111110110","000000000000001111","000000000000101100","111111111111110110","111111111111110110","000000000000001111","000000000000001001"),
("000000000000000001","111111111111111001","000000000000011101","000000000000010100","111111111111111000","111111111111101011","000000000000100000","111111111111011101","000000000000100110","111111111111101100","000000000000000011","111111111111101100","000000000000010001","000000000000110010","000000000000100011","000000000000000011","111111111111010110","000000000000011100","000000000000011010","000000000000001100","000000000000100001","111111111111111100","000000000000011100","111111111111101000","000000000000011000","111111111111101001","111111111111110101","000000000000100000","111111111111101110","000000000000000001","111111111111110110","000000000000100101","111111111111100111","000000000000000000","111111111111110110","111111111111010110","000000000000001011","111111111111110101","111111111111100101","000000000000001001","000000000000011011","000000000000010110","000000000000101101","000000000000010110","111111111111011100","000000000000001011","000000000000111010","111111111111100000","000000000000001010","000000000000100011","111111111111001001","111111111111011000","000000000000011011","111111111111111100","000000000000000110","000000000000000000","111111111111110010","000000000000011000","000000000000001101","000000000000010000","000000000000010010","000000000000000001","111111111111100101","111111111111110111","000000000000010110","000000000000110001","000000000000000111","111111111111011000","000000000000011010","000000000000001100","111111111111111101","000000000000101101","000000000000101011","000000000000010000","111111111111111111","111111111111111000","111111111111100010","000000000000000110","000000000000100001","111111111111110010","111111111111100010","111111111111101011","111111111111011110","000000000000110000","111111111111101011","000000000000000110","000000000000100011","000000000000000011","000000000000010001","111111111111111001","111111111111110011","111111111111111101","000000000000011110","111111111111111001","000000000000000111","111111111111110111","111111111111110011","000000000000001110","000000000000000010","000000000000100011","000000000000001001","111111111111101100","000000000000000110","111111111111011010","000000000000100101","111111111111010110","111111111111111111","000000000000010001","111111111111101001","000000000000010001","000000000000011101","111111111111111010","111111111111100011","000000000000010001","111111111111101000","000000000000101001","111111111111100110","000000000000011100","111111111111011011","111111111111111101","000000000000001111","111111111111111000","000000000000110101","000000000000010000","000000000000001100","111111111111011110","000000000000110011","111111111111110110"),
("111111111111111100","111111111111011101","000000000000011001","000000000000000111","111111111111010011","111111111111110100","000000000000011111","111111111111110011","000000000000000101","111111111111100101","000000000000010100","111111111111101101","000000000000011001","000000000000111110","000000000000010011","111111111111110111","111111111111011100","000000000000001111","000000000000000010","000000000000000100","000000000000101101","000000000000010001","000000000000101110","111111111111111110","000000000000011110","000000000000001101","111111111111010010","000000000000001111","000000000000000000","000000000000001100","111111111111111001","000000000000100010","000000000000001011","111111111111111100","000000000000010000","111111111111110111","000000000000001111","111111111111101101","000000000000001000","000000000000010000","000000000000010100","000000000000010110","000000000000010110","111111111111110111","000000000000001000","111111111111111011","000000000000000100","111111111111101001","000000000000000011","000000000000000010","111111111111001011","000000000000000110","000000000000000010","000000000000011000","000000000000000000","000000000000001111","000000000000010100","000000000000000100","000000000000001110","111111111111101100","000000000000001110","111111111111110000","111111111111111110","111111111111110101","000000000000100101","000000000000011100","000000000000010111","000000000000000101","000000000000001101","111111111111111110","000000000000000001","000000000000001010","000000000000011010","111111111111111101","000000000000001101","000000000000010011","000000000000000111","000000000000001000","000000000000000110","111111111111111101","111111111111110110","111111111111111111","111111111111101011","000000000000101111","111111111111111001","111111111111110001","000000000000000111","000000000000000100","000000000000010011","000000000000001101","111111111111011111","111111111111101111","000000000000110101","111111111111101111","000000000000010110","111111111111111000","000000000000000000","000000000000010011","000000000000001110","111111111111111100","111111111111111110","000000000000001001","000000000000001111","111111111111110000","111111111111110111","111111111111001111","000000000000000011","000000000000000000","000000000000000001","111111111111111011","111111111111111100","000000000000000100","111111111111110101","111111111111101111","111111111111111101","000000000000100001","111111111111101100","000000000000010100","000000000000001010","000000000000001011","000000000000001000","000000000000010000","000000000000001110","000000000000010111","111111111111101011","111111111111111100","000000000000010110","111111111111110010"),
("000000000000000001","111111111111001010","000000000000010001","000000000000000101","111111111111110111","111111111111110011","000000000000000011","111111111111100000","111111111111110101","111111111111110100","111111111111111000","111111111111101110","000000000000010000","000000000000011101","000000000000001001","000000000000011011","111111111111100010","000000000000000000","000000000000000100","111111111111101111","000000000000010100","000000000000000010","111111111111111001","000000000000001001","000000000000010111","111111111111111111","111111111111111100","000000000000011100","111111111111110001","000000000000001101","000000000000000010","000000000000010111","000000000000010010","111111111111110110","111111111111101101","111111111111101001","000000000000000100","111111111111111101","111111111111110111","000000000000000011","000000000000100100","111111111111101010","000000000000100011","000000000000001000","111111111111111000","111111111111100010","111111111111101000","111111111111110000","000000000000010010","000000000000001010","111111111111110000","111111111111110001","000000000000011001","000000000000100000","111111111111111011","000000000000010100","000000000000010001","111111111111111011","000000000000001100","111111111111111100","000000000000101110","111111111111110100","111111111111101111","000000000000010101","000000000000001101","000000000000101110","000000000000000110","111111111111110001","111111111111111101","000000000000000100","111111111111101111","000000000000001011","000000000000101010","111111111111111111","000000000000001010","111111111111110111","000000000000000001","111111111111110100","111111111111111111","111111111111101010","000000000000010000","000000000000000110","111111111111101110","000000000000000000","111111111111100110","000000000000010101","000000000000000111","111111111111101011","111111111111111111","000000000000000000","111111111111101100","111111111111110110","000000000000001101","111111111111111100","000000000000010101","111111111111110110","111111111111110101","000000000000011101","111111111111110110","111111111111111010","000000000000000001","000000000000000000","000000000000010100","111111111111101100","000000000000001001","111111111111100000","000000000000001010","000000000000010011","111111111111111011","000000000000011000","000000000000100000","111111111111101100","000000000000000010","111111111111101110","000000000000001000","000000000000010011","111111111111101100","111111111111111000","000000000000000111","000000000000010011","000000000000001001","000000000000001111","111111111111111011","000000000000100101","000000000000001000","000000000000000000","000000000000011011","000000000000010101"),
("000000000000000000","111111111111011001","000000000000001011","111111111111010011","111111111111001111","111111111111100101","000000000000100011","111111111111100110","000000000000011111","000000000000001110","000000000000011111","111111111111100101","000000000000010000","000000000000101111","000000000000001110","000000000000001011","111111111111010000","000000000000000011","000000000000100001","000000000000100001","000000000000010001","000000000000111101","000000000000101001","111111111111100101","000000000000001111","111111111111100101","111111111111110111","000000000000001101","000000000000000101","000000000000000101","111111111111111010","000000000000011110","111111111111110011","111111111111101011","000000000000010011","111111111111110101","000000000000101000","111111111111111000","111111111111101111","000000000000011110","000000000000111111","111111111111110101","000000000001000011","000000000000000111","111111111111100101","000000000000011001","000000000000010001","111111111111011110","000000000000010110","000000000000100110","111111111111101011","111111111111101001","000000000000011110","000000000000010100","000000000000000010","000000000000001100","111111111111011100","000000000000101000","000000000000001111","000000000000000001","000000000000001010","111111111111110101","111111111111101111","111111111111111011","111111111111011111","000000000000010110","000000000000000000","111111111111111111","111111111111111011","000000000000101111","111111111111011011","000000000000101011","111111111111110000","000000000000010111","111111111111111000","111111111111100001","111111111111101010","000000000000000110","000000000000001001","111111111111110001","111111111111011111","111111111111010100","111111111111101010","000000000000000001","111111111111110000","000000000000101000","000000000000100001","111111111111111001","111111111111110101","000000000000000100","111111111111111010","111111111111111100","000000000001000001","111111111111111100","000000000000100011","111111111111111111","111111111111111111","000000000000001000","000000000000001010","000000000000100111","000000000000000110","111111111111001010","111111111111101111","111111111111111100","000000000000011110","111111111111010011","111111111111110100","000000000000011101","111111111111010001","000000000000010011","000000000000011000","111111111111110111","111111111111010000","000000000000010011","000000000000001101","111111111111101111","111111111111100001","000000000000100011","111111111111100111","000000000000100010","000000000000001011","000000000000000110","000000000000011011","000000000000110110","000000000000001110","111111111111110101","000000000000100001","111111111111110011"),
("000000000000100011","111111111111101110","000000000000010001","111111111111111110","111111111111000011","111111111111100100","000000000000011001","111111111111100100","000000000000100000","111111111111111001","000000000000010100","111111111111010101","000000000000001101","000000000001001110","000000000000010001","111111111111110011","111111111111001011","000000000000011011","000000000000000100","000000000000001111","000000000001000000","000000000001011111","000000000000010010","111111111111110110","000000000000101110","000000000000001101","111111111111010111","111111111111111110","111111111111111001","111111111111101111","000000000000011011","000000000001000101","111111111111111101","000000000000001100","000000000000000100","111111111111111000","000000000000000000","111111111111010010","000000000000000100","111111111111100101","000000000000010011","111111111111111100","000000000000101011","000000000000111100","111111111111101001","111111111111011001","111111111111110111","111111111111001111","000000000000000011","000000000000100000","111111111110111110","111111111111001100","000000000000100011","000000000000110101","000000000000000101","000000000000001010","000000000000010100","000000000000101111","000000000000111111","000000000000001100","000000000000100100","111111111111110001","000000000000000111","000000000000000101","000000000000110110","000000000000101111","000000000000101111","111111111111111110","000000000000000100","111111111111100010","000000000000011000","000000000000010000","000000000000101000","000000000000110000","000000000000001011","000000000000001111","111111111111100110","000000000000100101","000000000000100000","111111111111101000","111111111111100110","111111111111101111","111111111111101000","111111111111101111","111111111111111011","111111111111110000","111111111111110100","111111111111001100","111111111111111010","111111111111011001","111111111111100011","111111111111111011","000000000001001110","111111111111110001","000000000000101010","000000000000110010","000000000000011101","000000000000111010","111111111111111011","000000000000010110","111111111111110100","111111111111111000","000000000000010111","111111111111111010","000000000000000110","111111111111001110","000000000000011100","000000000000101100","111111111111101110","000000000000000000","000000000000111110","111111111111000011","111111111111100001","111111111111110101","111111111111101011","000000000000000101","111111111111111101","000000000000001111","111111111111101110","000000000000111001","000000000000000110","111111111111111111","000000000000011110","000000000000001100","111111111111111001","000000000000001000","000000000000100101","000000000000001101"),
("000000000000100001","111111111111101010","000000000000011011","000000000000000000","111111111111001010","000000000000010000","111111111111111100","111111111111111101","000000000000011001","111111111111110111","111111111111110101","111111111111010011","000000000000000110","000000000000101101","000000000000000000","111111111111110100","111111111111011010","000000000000011011","000000000000001111","000000000000001001","000000000000010111","000000000000010010","000000000000101100","111111111111110111","000000000000011110","111111111111111110","111111111111100010","111111111111110110","111111111111101101","111111111111101000","000000000000010010","000000000000101000","000000000000000110","111111111111110101","111111111111110010","000000000000010100","000000000000001011","111111111111100001","000000000000010001","111111111111110110","111111111111111000","000000000000000100","000000000000001010","000000000000101011","000000000000000101","111111111111110001","000000000000011000","111111111111110110","111111111111111110","000000000000011001","111111111111110111","111111111111100101","000000000000010100","000000000000011000","000000000000000011","000000000000010100","000000000000000010","111111111111111011","000000000000001100","111111111111110111","000000000000110010","000000000000001101","111111111111101001","000000000000000100","000000000000010001","000000000000101110","000000000000010010","000000000000001011","000000000000100110","111111111111110001","000000000000001111","111111111111111011","000000000000100100","000000000000011110","000000000000010000","000000000000100111","111111111111111100","000000000000010010","111111111111111111","111111111111110011","000000000000001100","111111111111111000","111111111111111101","000000000000000000","111111111111100101","111111111111110010","000000000000000111","111111111111100010","000000000000010101","000000000000001011","111111111111001110","000000000000011101","000000000000000111","111111111111111010","000000000000010110","000000000000100011","000000000000011001","000000000000101001","111111111111111011","000000000000101010","111111111111111000","111111111111111010","000000000000000110","000000000000000101","000000000000000000","111111111111101100","000000000000010111","000000000000001100","000000000000011011","111111111111110111","000000000000011100","111111111111000110","000000000000000101","111111111111100101","111111111111111001","000000000000001110","000000000000010011","000000000000000000","000000000000010101","000000000000000111","000000000000001000","111111111111101011","000000000000100100","111111111111101101","111111111111100000","000000000000000110","000000000000100001","000000000000010110"),
("000000000000100111","111111111111101000","000000000000001100","000000000000010110","111111111111100101","111111111111111110","000000000000011011","111111111111010001","000000000000010010","111111111111111010","000000000000010100","111111111111010101","000000000000001000","000000000000010010","000000000000101111","111111111111110101","111111111111100110","000000000000101001","000000000000011011","111111111111111011","000000000000010000","000000000000000110","111111111111111100","111111111111110100","000000000000101000","000000000000000000","111111111111011000","111111111111101110","000000000000001010","000000000000011111","000000000000000001","000000000000011110","111111111111110011","111111111111111111","111111111111110101","000000000000000011","000000000000011001","111111111111001100","111111111111111101","000000000000000110","000000000000100111","000000000000010100","000000000000010000","000000000000001100","111111111111111001","000000000000000111","000000000000011011","111111111111100110","000000000000000100","000000000000110100","111111111111101101","111111111111011110","000000000000011000","000000000000100011","000000000000000111","000000000000000000","111111111111110101","000000000000001111","000000000000101000","000000000000000111","000000000000100110","111111111111111001","111111111111101010","111111111111100110","000000000000101001","000000000000011100","000000000000000001","111111111111111111","000000000000001001","000000000000001011","111111111111110101","000000000000000000","000000000000001001","000000000000010111","000000000000000111","000000000000010000","111111111111110111","111111111111101110","000000000000010111","000000000000000001","111111111111110000","111111111111011110","111111111111110010","000000000000100111","111111111111010001","000000000000001101","000000000000010100","111111111111011110","000000000000010000","000000000000001111","111111111111111101","111111111111111010","000000000000100001","000000000000000001","000000000000011100","000000000000000001","000000000000100001","000000000000011110","000000000000000001","000000000000100100","111111111111111111","111111111111111110","111111111111101001","111111111111101100","000000000000011001","111111111111010011","111111111111110110","000000000000101100","111111111111100010","000000000000001001","000000000000000110","111111111111100101","111111111111101101","000000000000010000","000000000000010000","000000000000000111","111111111111110110","000000000000010010","000000000000000011","000000000000010111","000000000000011111","111111111111101011","000000000000011101","000000000000001101","111111111111101011","000000000000000110","000000000000101101","111111111111110101"),
("000000000000100000","111111111111111000","000000000000010011","111111111111111110","111111111111101000","111111111111100001","000000000000100010","111111111111011010","000000000000001011","000000000000001010","111111111111101110","111111111111010000","000000000000000101","000000000000000000","000000000000101010","000000000000010010","111111111111101111","000000000000001101","000000000000000110","000000000000001101","000000000000011100","000000000000111110","000000000000100010","111111111111110010","000000000000010100","111111111111010001","111111111111110111","000000000000000000","000000000000000000","111111111111111001","111111111111100111","000000000000101110","111111111111101100","111111111111110100","111111111111110001","111111111111110011","000000000000101101","111111111111100111","111111111111110001","000000000000011101","000000000000110001","111111111111110110","000000000000110110","111111111111101110","111111111111110001","111111111111110000","111111111111101011","111111111111100000","000000000000001011","000000000000100000","111111111111101011","111111111111011000","000000000000010101","000000000000000100","000000000000011101","000000000000000000","111111111111111001","000000000000011101","000000000000100011","111111111111101110","000000000000000000","111111111111110001","000000000000001110","111111111111101111","000000000000000000","000000000000100100","000000000000010100","111111111111101010","000000000000011100","000000000000001110","111111111111100000","000000000000010101","111111111111101001","000000000000100101","111111111111111110","000000000000000000","111111111111111000","000000000000000001","000000000000100000","000000000000000000","111111111111011110","111111111111110101","111111111111100111","111111111111101100","111111111111010110","000000000000101100","000000000000101100","111111111111110000","111111111111111100","000000000000000011","000000000000001110","111111111111101010","000000000000100110","000000000000001001","000000000000011100","111111111111110100","111111111111110111","000000000000001001","000000000000000001","000000000000010111","111111111111101011","111111111111110000","111111111111110101","111111111111101101","111111111111111110","111111111111101111","111111111111111101","000000000000011110","111111111111111101","000000000000011011","000000000000011011","111111111111101110","111111111111001100","000000000000011011","000000000000010001","000000000000001010","111111111111101011","000000000000001011","111111111111100110","000000000000011010","000000000000001000","111111111111111011","000000000000100111","000000000001000010","000000000000000101","111111111111101111","000000000000000011","000000000000000001"),
("000000000000010100","000000000000001010","000000000000100101","000000000000010000","111111111111001100","111111111111111001","000000000000010001","111111111111000011","000000000000000000","000000000000000011","111111111111010100","111111111111100010","000000000000010001","000000000000100011","000000000000100101","111111111111110000","111111111111111001","111111111111110101","111111111111110011","000000000000010111","000000000000010001","000000000000001001","000000000000001001","000000000000000111","000000000000100010","111111111111111010","111111111111101011","000000000000000001","111111111111111100","000000000000010010","000000000000010101","000000000000011111","000000000000001000","111111111111110011","000000000000000000","111111111111110001","000000000000010100","111111111111111100","000000000000000000","111111111111111000","111111111111111011","111111111111101110","000000000000101001","000000000000100100","000000000000001011","000000000000000000","111111111111111101","111111111111011101","000000000000001110","000000000000011001","111111111111111100","000000000000000001","000000000000000101","000000000000100101","111111111111110110","000000000000001101","111111111111110101","000000000000100001","000000000000101011","000000000000001111","000000000000011101","111111111111101111","000000000000001010","111111111111111001","000000000000010101","000000000000101011","000000000000001100","111111111111101011","111111111111110001","111111111111101010","000000000000010011","111111111111101010","000000000000000000","000000000000011100","000000000000011000","111111111111111101","000000000000000110","000000000000010100","000000000000001100","000000000000000001","111111111111111111","000000000000001101","000000000000000011","111111111111100010","111111111111011100","000000000000100000","111111111111110010","111111111111101101","111111111111111111","111111111111010101","111111111111111110","111111111111110100","000000000000101000","111111111111111001","000000000000111010","111111111111110011","111111111111011111","000000000000001000","111111111111111000","000000000000001011","000000000000000010","000000000000000110","111111111111110111","000000000000001110","000000000000001110","111111111111000110","000000000000001001","111111111111111111","000000000000000000","000000000000011110","000000000000010100","000000000000000100","111111111111011100","000000000000000010","111111111111101101","111111111111111000","000000000000001101","111111111111111110","000000000000010001","000000000000000001","000000000000000000","111111111111111010","000000000000011110","000000000000011111","111111111111101111","000000000000000000","000000000000000001","111111111111111010"),
("000000000000000000","000000000000001101","000000000000011000","111111111111111011","111111111111010111","000000000000000000","000000000000101001","111111111111010011","111111111111111110","111111111111111100","111111111111100110","111111111111100110","000000000000000100","000000000000000001","000000000000000100","111111111111011011","111111111111110001","111111111111101100","000000000000001100","000000000000001111","000000000000001011","000000000000001010","111111111111110111","000000000000000000","000000000000101000","111111111111110011","111111111111100010","000000000000010101","111111111111101000","111111111111110001","000000000000011000","000000000000101010","111111111111111011","111111111111111001","111111111111111111","000000000000000011","000000000000001000","111111111111110110","000000000000010111","111111111111101111","000000000000010101","111111111111110010","000000000000000000","000000000000010011","111111111111101001","111111111111110110","111111111111101011","111111111111100011","111111111111101000","000000000000011000","111111111111110000","111111111111110100","000000000000000110","000000000000001010","000000000000000111","000000000000010101","000000000000000000","000000000000001000","000000000000110010","000000000000001110","000000000000001011","111111111111110011","000000000000001100","000000000000001111","000000000000001010","000000000000001010","000000000000000110","111111111111110100","111111111111100011","111111111111101100","111111111111111000","111111111111111000","111111111111110011","000000000000011111","000000000000000011","111111111111110111","000000000000000101","000000000000001000","000000000000001110","111111111111111101","000000000000010001","000000000000010000","111111111111110110","111111111111011011","111111111111010110","000000000000001100","111111111111111011","111111111111110110","000000000000001111","111111111111100110","111111111111110000","000000000000010100","000000000000110001","000000000000010010","000000000000110100","111111111111111000","111111111111101010","000000000000011010","111111111111110110","111111111111111100","111111111111110101","111111111111100110","111111111111110000","111111111111101110","000000000000010101","111111111111101111","000000000000100010","111111111111111101","000000000000010000","000000000000011001","000000000000110100","000000000000001001","111111111111011110","111111111111100010","111111111111101101","111111111111111100","000000000000000001","000000000000001100","111111111111110111","000000000000000001","111111111111111001","111111111111111111","000000000000010101","000000000000010011","111111111111100101","000000000000010101","111111111111111110","000000000000011000"),
("111111111111110111","000000000000000101","111111111111111001","000000000000000101","000000000000001000","000000000000000010","000000000000010101","000000000000000000","111111111111101110","000000000000001100","111111111111100000","111111111111110000","000000000000011111","000000000000010110","000000000000000110","000000000000000000","000000000000000000","111111111111101010","111111111111101111","000000000000000000","000000000000010110","000000000000011101","000000000000011010","111111111111110010","111111111111111000","111111111111110011","000000000000001110","000000000000001101","111111111111111110","000000000000000110","111111111111100110","000000000000000000","000000000000001110","000000000000000111","111111111111110010","111111111111111111","000000000000011101","111111111111111000","000000000000000101","000000000000000101","000000000000000000","000000000000000100","111111111111110101","000000000000011101","111111111111111110","000000000000000101","111111111111101100","111111111111110100","000000000000010011","111111111111111110","111111111111101111","111111111111111101","111111111111111000","000000000000001110","000000000000010100","000000000000001001","111111111111101111","000000000000001011","000000000000011001","111111111111111010","111111111111110111","000000000000001101","000000000000000111","000000000000000111","111111111111110100","000000000000000011","000000000000010000","111111111111111000","111111111111100000","000000000000011010","111111111111101101","000000000000000100","111111111111100101","000000000000011011","111111111111111001","111111111111111111","111111111111110011","000000000000010010","000000000000010011","000000000000001100","111111111111110101","000000000000000100","000000000000000011","000000000000001001","111111111111101111","111111111111111000","111111111111111100","000000000000000100","000000000000000000","000000000000000110","111111111111110101","111111111111011111","111111111111101010","000000000000000010","000000000000010100","000000000000001000","111111111111101010","111111111111110011","000000000000010000","111111111111110101","111111111111100011","000000000000000001","000000000000001100","111111111111101101","000000000000000000","000000000000000000","000000000000000100","111111111111110001","111111111111110000","000000000000001000","111111111111111111","000000000000000000","111111111111111000","111111111111111110","111111111111111110","111111111111110110","000000000000000111","111111111111110111","000000000000000101","111111111111111100","111111111111111111","111111111111111110","000000000000100001","000000000000001100","111111111111111101","111111111111101111","111111111111111111","111111111111101101"),
("000000000000000101","111111111111101000","000000000000001010","000000000000010110","000000000000000111","111111111111111010","000000000000011101","111111111111111111","111111111111110011","000000000000011001","111111111111001101","111111111111010011","000000000000011010","000000000000000101","000000000000100101","000000000000000010","000000000000000110","111111111111111101","111111111111110100","111111111111110100","000000000000010100","000000000000101000","000000000000000000","111111111111111010","111111111111101000","111111111111111111","111111111111011111","111111111111111011","111111111111111010","111111111111110011","111111111111101101","000000000000100100","111111111111110010","111111111111010001","000000000000000000","111111111111110010","000000000000010000","111111111111100111","111111111111011001","111111111111111101","000000000000011010","000000000000010000","000000000000100010","000000000000001110","111111111111101000","111111111111111110","111111111111100011","111111111111100100","000000000000000101","111111111111110111","000000000000011001","111111111111101000","000000000000100110","111111111111110001","111111111111100111","000000000000101101","111111111111111111","000000000000001111","000000000000101110","000000000000001001","111111111111110011","111111111111101111","111111111111110000","111111111111101100","111111111111101111","000000000000010001","000000000000010010","111111111111111000","000000000000010111","000000000000100000","111111111111100001","111111111111111101","111111111111110100","000000000000010001","111111111111101010","111111111111010100","111111111111100000","111111111111110101","000000000000011100","111111111111110101","111111111111100101","111111111111110010","111111111111101010","000000000000000001","000000000000000000","000000000000100111","000000000000100000","111111111111110011","111111111111101001","111111111111101111","000000000000011000","111111111111010111","111111111111010101","000000000000000001","000000000000010001","000000000000000000","111111111111111100","111111111111110100","111111111111111010","000000000000100001","111111111111110111","111111111111011001","000000000000010000","111111111111110111","000000000000010001","111111111111100011","000000000000010111","000000000000000101","000000000000001111","000000000000100110","000000000000011111","111111111111100111","111111111111100011","000000000000010110","000000000000000000","000000000000001100","111111111111111100","000000000000001110","111111111111110000","000000000000001100","111111111111110011","111111111111101010","111111111111111110","000000000000010101","000000000000100111","111111111111110111","000000000000000111","111111111111100101"),
("111111111111110000","111111111111101101","111111111111111011","000000000000011101","111111111111110010","111111111111111100","000000000000010101","000000000000010000","000000000000000111","000000000000101010","111111111111011000","111111111111011010","000000000000001001","000000000000001100","000000000000011000","111111111111101010","111111111111110000","000000000000000100","111111111111011010","000000000000001110","000000000000010001","000000000000101110","111111111111100010","111111111111111101","111111111111011111","111111111111101000","000000000000000001","000000000000001011","000000000000001101","111111111111111000","111111111111110110","000000000000101000","000000000000001111","111111111111010110","000000000000010011","000000000000000100","000000000000011101","111111111111100101","111111111111111001","000000000000001001","000000000000011100","000000000000011111","000000000000010110","000000000000111000","111111111111101010","000000000000001011","111111111111010100","111111111111101011","000000000000001101","111111111111111011","000000000000101110","111111111111110000","000000000000100111","000000000000001000","111111111111100000","000000000000001101","111111111111100011","000000000000000100","000000000000011100","000000000000001000","111111111111110001","000000000000000110","111111111111101010","111111111111110011","111111111111110001","000000000000001101","000000000000010011","111111111111100110","000000000000001101","000000000000010000","111111111111101011","111111111111100110","111111111111100111","000000000000101100","111111111111110000","111111111111010000","111111111111110111","000000000000001010","000000000000100100","000000000000011111","111111111111111111","111111111111011011","111111111111111010","111111111111110010","000000000000000111","000000000000100100","000000000000001011","111111111111101101","111111111111101110","000000000000001100","000000000000011000","111111111111101100","111111111111110011","111111111111110000","000000000000010010","000000000000010001","111111111111110101","111111111111111100","000000000000010001","000000000000011011","111111111111011100","111111111111100010","000000000000001000","000000000000000000","000000000000011110","111111111111111101","111111111111110011","111111111111110000","111111111111110000","000000000000110011","000000000000100100","000000000000000000","111111111111111101","000000000000011000","000000000000100000","000000000000000111","111111111111111010","000000000000000010","000000000000000011","111111111111110100","111111111111110010","111111111111110110","000000000000000100","000000000000100011","000000000000001101","111111111111100000","111111111111101010","000000000000000010"),
("000000000000001010","111111111111111010","000000000000011011","000000000000001100","000000000000011001","111111111111011111","111111111111111011","111111111111110011","111111111111111111","000000000000011110","000000000000000111","111111111111100100","000000000000000101","000000000000011001","000000000000100101","000000000000001111","000000000000000110","000000000000100101","000000000000001001","111111111111111000","000000000000001100","000000000000101011","000000000000001111","000000000000001111","111111111111011011","111111111111011100","000000000000000001","000000000000010010","000000000000000111","000000000000010000","111111111111101011","111111111111111011","111111111111110110","000000000000001111","000000000000011000","111111111111110111","000000000000100000","111111111111111101","000000000000000100","000000000000100010","000000000000011111","000000000000000101","000000000000000110","000000000000000111","111111111111011101","111111111111101101","111111111111110001","111111111111111101","000000000000100101","000000000000011000","000000000000100101","000000000000000010","000000000000010100","111111111111100100","111111111111110010","000000000000100010","111111111111111011","111111111111111001","111111111111111100","000000000000000000","111111111111111100","000000000000000110","111111111111110000","111111111111100000","000000000000010011","000000000000000111","000000000000000000","000000000000001100","000000000000000101","000000000000011110","111111111111011011","000000000000010011","000000000000001000","000000000000000101","111111111111110000","111111111111101011","111111111111011010","111111111111110001","000000000000000100","000000000000010010","111111111111101110","111111111111011110","111111111111101100","000000000000000000","000000000000000001","000000000000011001","000000000000010011","111111111111110101","000000000000000110","111111111111111111","111111111111111110","111111111111111100","000000000000011110","111111111111111010","000000000000000111","111111111111110100","000000000000001100","000000000000010010","111111111111110000","000000000000011111","111111111111011101","111111111111111010","000000000000010001","111111111111110001","111111111111111100","111111111111101110","111111111111101111","000000000000000001","111111111111110100","000000000000001011","000000000000011101","111111111111110000","111111111111110111","000000000000000110","000000000000100111","111111111111100110","000000000000010001","111111111111111001","000000000000000110","000000000000000100","000000000000010001","111111111111100000","000000000000001010","000000000000001101","111111111111111010","111111111111111100","000000000000010110","111111111111011111"),
("111111111111111100","000000000000001000","000000000000010010","000000000000000000","000000000000000000","111111111111110011","111111111111110010","111111111111101111","000000000000000000","111111111111111100","000000000000001100","000000000000010100","111111111111110100","111111111111110110","000000000000001110","111111111111110010","000000000000000111","111111111111110101","000000000000000011","111111111111111000","111111111111111001","111111111111110000","000000000000001100","111111111111111010","111111111111110111","111111111111110111","111111111111110101","111111111111111001","000000000000001100","111111111111110000","000000000000010001","111111111111111001","111111111111110100","111111111111110100","000000000000000111","111111111111110011","000000000000001100","000000000000001011","111111111111111111","000000000000010000","111111111111101101","000000000000000001","111111111111110000","000000000000001111","111111111111110011","000000000000000100","000000000000000001","111111111111110101","111111111111111111","000000000000001100","000000000000001101","111111111111111000","111111111111110000","111111111111110101","000000000000000001","000000000000000100","000000000000010100","000000000000001110","000000000000000000","000000000000000100","000000000000000000","000000000000001011","000000000000000010","000000000000010001","000000000000001100","111111111111110011","111111111111110010","000000000000001010","111111111111110010","000000000000000010","111111111111111000","000000000000000000","111111111111111001","111111111111111000","111111111111110111","111111111111101110","000000000000000000","000000000000010000","111111111111111101","000000000000000011","000000000000010100","111111111111111010","111111111111101111","111111111111111010","111111111111101110","000000000000010000","111111111111101101","000000000000001101","000000000000000000","111111111111110111","111111111111101111","000000000000001100","000000000000001111","000000000000001101","111111111111110011","111111111111111001","000000000000001101","111111111111111110","000000000000001101","000000000000001011","000000000000010001","000000000000001001","111111111111101111","000000000000000000","000000000000000000","000000000000000111","000000000000000011","111111111111111011","000000000000000010","111111111111110100","000000000000010000","111111111111110101","000000000000000111","000000000000000101","111111111111111111","111111111111110000","111111111111111100","000000000000001100","000000000000000110","000000000000001100","111111111111110111","000000000000010001","000000000000001010","000000000000000001","000000000000010000","111111111111101101","000000000000010010","000000000000010100"),
("000000000000000110","111111111111101101","000000000000000101","111111111111110000","000000000000010000","111111111111110110","000000000000000000","111111111111111100","000000000000000001","111111111111110011","000000000000000101","111111111111111111","000000000000000000","000000000000000001","111111111111110001","000000000000000011","111111111111110110","111111111111111110","111111111111111000","000000000000000001","111111111111110000","000000000000001011","000000000000001111","000000000000000110","111111111111111100","111111111111101110","000000000000001100","000000000000010010","000000000000001011","111111111111111111","111111111111110011","000000000000000111","111111111111110100","111111111111110001","111111111111110010","111111111111110010","111111111111111110","000000000000000111","111111111111111001","111111111111111000","000000000000001100","000000000000000000","111111111111110110","111111111111101101","111111111111111101","000000000000001110","111111111111111110","111111111111111010","000000000000000000","000000000000000010","111111111111110101","111111111111111101","000000000000010001","111111111111101111","111111111111101101","000000000000000100","000000000000001101","000000000000000101","000000000000000110","111111111111110101","000000000000001010","000000000000001111","111111111111111000","000000000000010011","000000000000001011","000000000000000000","111111111111110110","111111111111110000","111111111111111111","111111111111111111","000000000000001000","111111111111110000","000000000000000100","000000000000001000","111111111111111111","111111111111111101","111111111111101110","000000000000010010","000000000000000111","000000000000000011","111111111111110000","000000000000000000","000000000000000000","000000000000000001","000000000000001001","111111111111101101","111111111111101100","111111111111110101","000000000000000000","111111111111101101","000000000000000001","000000000000000111","000000000000000011","111111111111111001","000000000000010100","111111111111111000","000000000000000011","000000000000000011","111111111111101111","111111111111111001","111111111111110110","111111111111111101","000000000000000101","000000000000000110","111111111111110110","000000000000010011","000000000000010010","111111111111110010","111111111111110011","000000000000001101","111111111111101110","000000000000001000","000000000000000000","111111111111101110","111111111111110101","000000000000000010","111111111111111101","000000000000010010","111111111111111110","000000000000000010","111111111111111000","111111111111101100","111111111111110111","111111111111111101","111111111111111000","000000000000000000","111111111111111101","111111111111110101"),
("000000000000010011","000000000000001101","111111111111111111","111111111111110000","111111111111101111","000000000000000011","111111111111110001","000000000000001011","000000000000001000","000000000000010000","000000000000000111","111111111111111011","111111111111110110","111111111111101110","000000000000001110","000000000000001011","000000000000001111","000000000000001111","111111111111110100","000000000000010011","000000000000000100","000000000000000111","111111111111101110","111111111111111111","111111111111111101","000000000000010001","111111111111111010","111111111111111000","111111111111111000","000000000000000011","000000000000001011","000000000000001110","000000000000001001","000000000000000110","111111111111101100","000000000000001000","111111111111110111","111111111111111000","111111111111110110","111111111111111001","111111111111111100","111111111111111101","111111111111110100","111111111111111110","000000000000001110","000000000000010001","000000000000000000","000000000000000101","111111111111111111","111111111111111000","000000000000000010","000000000000001010","000000000000000010","000000000000010001","111111111111111010","111111111111111111","000000000000000001","111111111111101101","111111111111110011","000000000000001110","000000000000001010","000000000000010010","000000000000000000","000000000000000011","000000000000001011","111111111111110100","000000000000000110","000000000000000101","111111111111101110","111111111111110111","111111111111110101","000000000000010001","111111111111101100","000000000000010000","111111111111111100","000000000000001110","000000000000000100","000000000000010011","111111111111101101","000000000000000000","000000000000001000","111111111111101100","000000000000001011","000000000000010011","000000000000000100","000000000000001010","111111111111110100","111111111111111010","000000000000010001","111111111111101111","111111111111111000","111111111111110000","000000000000000111","000000000000001110","111111111111111111","000000000000010011","000000000000001011","111111111111110101","111111111111110101","111111111111110010","111111111111110100","111111111111110100","000000000000010100","111111111111111111","111111111111110100","000000000000010001","000000000000010010","111111111111101111","111111111111111001","111111111111111110","000000000000001000","111111111111111001","000000000000000011","000000000000000010","111111111111111101","111111111111111110","111111111111101111","111111111111101110","000000000000000001","000000000000001011","000000000000001001","000000000000000011","000000000000001100","111111111111110010","000000000000010100","111111111111111010","000000000000001010","111111111111110011"),
("000000000000001011","111111111111111100","111111111111110010","111111111111111010","000000000000010010","111111111111111110","000000000000000001","111111111111101110","000000000000000011","111111111111111110","111111111111110001","000000000000000100","111111111111111101","000000000000001110","000000000000010010","000000000000001111","111111111111101111","000000000000000110","111111111111111001","000000000000010010","111111111111111011","111111111111111000","000000000000001010","111111111111111110","000000000000000001","111111111111101100","111111111111111111","000000000000000000","000000000000001110","111111111111110001","000000000000001000","111111111111111100","111111111111101110","000000000000010000","111111111111101100","111111111111101110","000000000000010000","000000000000001111","111111111111110011","111111111111110010","000000000000000000","000000000000000001","111111111111101110","111111111111110111","111111111111110110","111111111111110111","000000000000001011","111111111111110110","000000000000010001","000000000000001100","000000000000000001","111111111111110000","000000000000001000","111111111111110001","111111111111111101","000000000000001101","000000000000000010","000000000000001110","111111111111111011","000000000000000110","000000000000001111","111111111111111000","000000000000001010","111111111111101100","000000000000010001","111111111111110001","000000000000001000","000000000000001010","111111111111110100","000000000000001011","000000000000000000","000000000000010001","111111111111111101","111111111111110011","111111111111110011","000000000000001101","000000000000010010","000000000000000001","000000000000001011","111111111111111010","111111111111110010","111111111111110000","000000000000010011","111111111111111110","111111111111101101","000000000000000101","111111111111110100","000000000000000100","000000000000001101","111111111111111000","000000000000010100","000000000000000111","111111111111101101","000000000000000000","111111111111110010","000000000000000100","111111111111110100","000000000000010000","111111111111101110","111111111111110000","111111111111111011","111111111111110000","000000000000001010","000000000000000011","111111111111110101","000000000000001100","111111111111110000","111111111111110010","111111111111111100","000000000000001110","111111111111111110","111111111111111111","000000000000000001","111111111111110011","111111111111111100","111111111111101111","000000000000001101","000000000000000110","111111111111110110","111111111111110000","000000000000010010","111111111111111111","111111111111110110","111111111111111111","000000000000000010","000000000000000111","000000000000010100","000000000000000100"));

	constant weights_2 : weight_2 := (("111111111101110001","111111111111101111","000000000000101010","111111111110000100","111111111111011100","000000000001000000","000000000001011001","111111111110001111","111111111111110110","000000000001000110"),
("000000000001010010","111111111111001100","111111111101000110","000000000000010000","000000000000111011","000000000000010101","000000000001001001","111111111111111110","111111111101111110","000000000001010000"),
("111111111110110000","111111111111100101","111111111111001010","111111111111111100","000000000000111101","000000000001010000","111111111101011101","000000000000111000","111111111111001111","000000000001000000"),
("111111111111111101","000000000000100110","000000000000111011","000000000000000111","111111111110010011","111111111111001101","111111111111010110","111111111111011001","000000000000100011","111111111111111000"),
("111111111111010011","000000000001100101","111111111101111001","111111111110011001","000000000010011100","111111111111011100","000000000000101011","111111111111011011","111111111111001101","111111111110000000"),
("111111111111000110","000000000000101000","000000000000101011","111111111111101110","000000000000101111","111111111111101100","000000000000111011","111111111110100100","000000000000010000","111111111111101110"),
("000000000000110011","111111111110111011","000000000000110100","111111111111001010","111111111111111110","111111111111001111","000000000000010111","000000000000011010","000000000000110000","000000000000110100"),
("000000000000001110","111111111111110110","000000000000001100","000000000000101010","000000000000001000","000000000000000100","111111111111010111","111111111110010001","000000000001100001","111111111111100110"),
("111111111110110001","000000000000010100","000000000000011111","000000000000011010","000000000000000101","111111111111001001","111111111110111100","000000000000011110","000000000000101010","000000000000010001"),
("000000000001000001","111111111111110101","111111111111101111","000000000001000111","111111111111111000","111111111111011100","000000000000010110","000000000001100001","111111111110011100","111111111110100000"),
("111111111111100001","000000000001010011","000000000001111110","000000000000100100","111111111111011011","000000000000001000","111111111111111001","000000000000000000","000000000000001001","111111111101011100"),
("000000000001000010","111111111111010011","111111111110111110","000000000000010100","111111111111001111","000000000001010101","000000000000100000","111111111111000101","000000000000101111","111111111111001001"),
("111111111111010010","000000000000111000","000000000000110111","000000000000001100","111111111110100000","000000000000000001","111111111110100110","000000000000100110","111111111111111100","000000000000100010"),
("111111111111111101","000000000001011110","111111111111000001","111111111111100100","111111111111001011","000000000001000011","111111111111000010","000000000000101001","111111111101101011","000000000001100000"),
("111111111110111001","111111111111001111","000000000000001010","111111111110010110","000000000000110001","111111111110001100","000000000001010110","000000000001001011","111111111111100110","000000000000011110"),
("000000000000011101","111111111111100011","000000000000111101","111111111111100111","111111111110010110","111111111111111111","000000000000001001","111111111111111010","111111111111011010","111111111110010101"),
("000000000000001110","000000000000000001","000000000000101111","000000000000101101","000000000000111011","111111111111001001","000000000000010111","111111111111100101","111111111111010110","111111111110011000"),
("000000000000000100","000000000000100001","000000000000101011","111111111111101010","111111111110010100","000000000000000000","111111111111010110","000000000000010001","000000000000101100","111111111111001100"),
("111111111110010010","111111111111111001","000000000000010010","111111111111111111","111111111110111100","111111111111101101","111111111111100001","000000000000110111","000000000000100101","111111111110100111"),
("000000000000010011","111111111111001101","000000000000110000","000000000000101001","000000000000011011","000000000000000011","111111111111001011","000000000000011111","111111111111001110","111111111110111100"),
("111111111111110110","000000000000011110","000000000000001111","111111111111010101","111111111101111101","000000000001000000","111111111101001101","000000000000110111","111111111111110111","000000000000100000"),
("000000000001000010","000000000001001111","000000000000000000","111111111110100011","000000000000001100","111111111111011001","111111111111001011","000000000010011111","111111111111100111","000000000000000110"),
("000000000001001101","000000000001101011","111111111111111111","111111111111110001","000000000001110010","111111111110100101","111111111111111100","000000000000101001","111111111110010100","111111111111110011"),
("000000000000101000","000000000000100001","111111111110101111","111111111101110000","000000000001000000","111111111111011010","111111111111011001","000000000000000111","000000000001000000","000000000000000111"),
("000000000000110101","111111111111000101","111111111111100010","111111111111000100","111111111111100111","000000000000110111","111111111111110011","000000000000001111","000000000000001110","000000000000011000"),
("111111111111001001","000000000000010100","000000000000101100","000000000000010000","111111111111111000","111111111111111001","000000000000010100","111111111111010001","000000000000101000","000000000000000111"),
("111111111110111011","000000000001000111","111111111111101001","111111111111011101","000000000001011001","000000000000100100","111111111110111000","111111111111011011","000000000000000101","111111111110001100"),
("000000000000011000","111111111111101011","000000000000111101","000000000000100111","111111111101111010","111111111111011000","111111111111100100","000000000000001110","111111111111110010","000000000000110111"),
("111111111110011010","000000000000110100","000000000000011110","000000000000110001","000000000000110111","111111111110001011","000000000000110011","000000000000110100","000000000000000011","111111111111001110"),
("000000000000111010","000000000000011101","111111111110110001","000000000000010000","111111111110100000","000000000001011001","000000000001001101","111111111111101101","111111111110110101","111111111110001100"),
("111111111111000000","000000000000011110","000000000000110011","111111111111111100","111111111111111110","000000000000111001","111111111111110110","111111111111011011","000000000000010110","000000000000101001"),
("111111111111010111","000000000000011000","111111111111001101","000000000000110101","111111111111001011","111111111111111100","000000000001010101","000000000000000110","111111111111011001","000000000000010100"),
("000000000000101100","111111111110111000","000000000000101101","000000000000110100","000000000000000110","000000000000101001","111111111111111010","000000000000000100","000000000000011011","000000000000100011"),
("000000000000101101","000000000001010000","111111111110100111","111111111111011110","111111111110111001","000000000001011010","000000000001100001","111111111111011000","000000000000000101","000000000000100111"),
("111111111111011001","000000000000100111","000000000000110100","111111111111010110","000000000000100100","000000000000101001","000000000000010110","000000000000101011","000000000000101011","111111111111101111"),
("111111111110000001","000000000000110010","111111111111011001","000000000000110001","000000000000101100","111111111111001001","111111111111000010","111111111110011011","000000000000111111","000000000000001110"),
("111111111111111100","111111111110110100","000000000000001010","111111111111010111","111111111111111000","000000000000110101","111111111111111100","000000000000110111","111111111111101011","000000000000000110"),
("111111111110111010","000000000000111010","000000000000011101","000000000000110000","000000000000111100","000000000000110101","111111111111001010","111111111111111001","000000000000100111","111111111111001010"),
("111111111110101011","000000000000101100","111111111110000111","000000000000010000","000000000001000000","000000000000101111","000000000000000101","111111111111011001","111111111111011111","000000000000100111"),
("111111111111100010","111111111111011110","111111111111011110","000000000000111000","000000000000100101","000000000000111000","111111111111010111","000000000000101110","111111111111011110","111111111111100111"),
("000000000000100010","000000000001011001","111111111111001100","000000000000000100","111111111110110011","000000000001001100","111111111111001000","000000000000100000","111111111110101010","111111111111101000"),
("111111111110000000","000000000000110100","111111111111101100","111111111110110000","000000000000011100","000000000000110111","000000000000101001","000000000000111101","000000000000100010","111111111111001101"),
("000000000010001010","000000000000011001","000000000001010111","111111111111100111","111111111110111100","111111111101000010","000000000001000111","000000000000110010","111111111111110101","000000000000010001"),
("000000000001000101","000000000000110100","000000000000110111","111111111111100010","111111111111110101","111111111110001110","000000000000111101","111111111111111001","000000000000000110","000000000000010110"),
("111111111111011010","111111111110110111","111111111111111010","000000000000010100","000000000000110000","000000000000010000","111111111111111100","111111111110111010","000000000000100100","000000000000000111"),
("111111111111010011","000000000001001011","111111111111100010","000000000000011001","000000000001010000","111111111111100110","000000000000011101","000000000000111110","111111111110010110","111111111111100110"),
("000000000000101101","000000000000010010","000000000000011110","000000000000001010","111111111111001100","111111111111010100","000000000001000100","000000000000110101","000000000000101000","111111111101001101"),
("111111111110101100","000000000001001000","000000000000110101","111111111110101000","000000000000000100","000000000000110101","000000000000110011","111111111111011110","000000000000111111","111111111110000010"),
("000000000000000001","111111111110110010","111111111111000111","000000000000011101","000000000000011100","000000000000101010","111111111111100100","000000000000101100","000000000000100010","111111111111101001"),
("111111111111110000","111111111111001110","111111111111000110","000000000000010100","111111111111110101","111111111110111010","000000000000101010","000000000000010110","000000000000001000","000000000000001001"),
("000000000000110001","000000000000010100","000000000000010100","000000000000011000","111111111111010010","111111111111001111","111111111111011110","111111111111110110","000000000001100100","111111111101110011"),
("000000000000101100","111111111111100100","000000000000101001","000000000000011110","000000000000110110","000000000000100000","111111111111101001","111111111111011001","000000000000100101","111111111111110001"),
("000000000000100101","111111111111001101","111111111111011010","111111111110110101","111111111111000101","111111111111110111","111111111111101101","000000000000101011","000000000000011011","111111111111100100"),
("111111111111010100","000000000000101100","111111111111111100","000000000000101101","111111111111000110","000000000000101110","111111111110011110","000000000000010011","000000000000000110","000000000001001011"),
("111111111111001100","000000000000100010","000000000000100010","000000000000111111","000000000000010000","000000000000101001","111111111101100111","000000000000111000","111111111111100010","000000000000101101"),
("111111111111001000","000000000000010101","000000000000110011","000000000000000010","000000000000111111","111111111111100010","111111111111001000","000000000000101101","000000000000100000","000000000000110011"),
("111111111111101100","111111111111111100","111111111110001000","000000000000010010","000000000000011000","000000000001000100","000000000000001111","000000000000000100","000000000000110011","000000000001000000"),
("000000000000011100","111111111110110010","000000000000000001","000000000000101010","111111111110111011","111111111111010101","111111111110110101","000000000000011011","111111111111100101","000000000000000011"),
("000000000000110001","111111111110110101","111111111111001101","111111111111100000","111111111111110011","111111111111001011","111111111111010000","000000000000010100","111111111111111111","000000000000010000"),
("000000000000000000","000000000000101010","000000000000010000","111111111111100000","111111111111111010","111111111111001110","000000000000011101","000000000000101011","000000000000100110","111111111111010010"),
("000000000000010001","111111111111011100","111111111111010110","000000000000100101","111111111110110100","000000000000001110","111111111111110000","111111111111111100","000000000000010101","000000000000011100"),
("111111111111110010","000000000000111011","000000000001101110","000000000001011101","111111111110010110","000000000000101110","111111111101111110","000000000001100100","111111111101111011","111111111110111011"),
("000000000000100101","000000000000011111","000000000001000110","000000000000010000","000000000000001000","111111111110111001","111111111110100111","000000000001011011","111111111111111010","111111111111000011"),
("000000000000010001","000000000001000001","111111111111111110","111111111111101101","000000000000101100","111111111110111110","000000000000001111","111111111111001000","000000000000100000","000000000000001111"),
("000000000000000100","000000000000111111","111111111110010110","111111111110011001","000000000000111001","111111111110010011","111111111110100001","111111111111011101","111111111110011110","000000000001110111"),
("000000000000110100","111111111110010111","111111111111011110","111111111111000111","000000000000011101","000000000000100110","000000000000000111","000000000000101001","000000000000100001","000000000000101110"),
("000000000000011000","111111111111010110","111111111101100011","111111111111010011","111111111110101001","000000000001100011","111111111111011101","111111111111011010","000000000000001001","111111111111111001"),
("000000000000000100","111111111111101001","000000000000000001","000000000000001010","111111111111011100","000000000000000000","000000000001000010","111111111110010111","000000000000011010","111111111111100010"),
("111111111110100110","111111111101110010","000000000000001101","000000000010101111","111111111110010000","000000000000110010","111111111101111001","000000000001010111","111111111110010001","111111111111001111"),
("000000000000011011","000000000000001000","111111111111111100","111111111111001101","000000000000110100","000000000001000100","111111111111111000","000000000001010111","111111111111110111","111111111110000000"),
("111111111111010101","000000000000100111","000000000000010000","000000000000100100","111111111111011110","111111111111011011","000000000000001111","111111111110111000","000000000000101101","000000000000001000"),
("111111111111101101","000000000000110000","000000000000001100","000000000000101001","111111111110011010","000000000000000011","111111111111010001","000000000000011001","000000000000001010","111111111111001111"),
("000000000000001011","111111111111110011","111111111111000100","000000000001000101","111111111101111111","000000000001111000","000000000000111110","111111111111100010","111111111111010001","000000000000011100"),
("000000000001001000","000000000000010000","000000000000100000","000000000000111001","111111111111110100","111111111110001001","111111111110001111","000000000000111001","111111111111110101","000000000000110000"),
("111111111101110100","000000000000100101","111111111111001111","000000000000011100","111111111111010000","000000000000001110","000000000000001011","111111111111100010","000000000000001011","000000000000001101"),
("111111111110111100","111111111110100110","000000000001001110","000000000001010010","111111111111011111","000000000000100100","000000000000010110","111111111110110011","111111111110010011","000000000000110101"),
("111111111111010101","111111111110111110","000000000000101010","111111111111001001","000000000000100111","000000000000100111","000000000000000101","111111111111100011","000000000000100011","000000000000001101"),
("000000000000010010","111111111111011110","000000000000111101","000000000000110111","111111111110001110","000000000000000101","111111111111000000","111111111111110010","111111111111101011","000000000000111001"),
("111111111111110111","111111111111000001","000000000000000111","111111111111010001","000000000000110101","111111111110111101","000000000000010000","000000000001000010","111111111111111001","000000000000100001"),
("000000000000010011","111111111111001111","000000000000100010","000000000000010000","000000000000110100","111111111111001011","000000000000000000","000000000000010100","000000000000010100","111111111111010101"),
("000000000000011000","000000000000110111","111111111110111010","111111111111001000","000000000000111001","000000000000011111","000000000000010111","111111111110111011","000000000000000111","000000000000001110"),
("000000000000001000","111111111110111011","000000000000001101","000000000000011000","000000000000010101","000000000000011101","111111111111111111","111111111111011000","000000000000011011","000000000000101101"),
("000000000000001111","000000000000100010","000000000001110110","111111111111110001","000000000001000110","111111111110111111","000000000000100001","111111111110111010","111111111110001100","000000000000010101"),
("111111111111100000","000000000001100010","111111111110101011","000000000000000110","000000000001000010","111111111111000000","111111111111101100","000000000001011110","111111111101110111","111111111101010110"),
("000000000000011111","000000000001000100","000000000000001100","000000000000101000","111111111111000111","000000000000000101","111111111111010101","111111111110101011","000000000000010110","111111111111011101"),
("000000000001000011","111111111111111101","000000000000001101","111111111111100101","000000000000110000","111111111111111001","000000000000010011","000000000000101000","111111111110010011","000000000000011011"),
("111111111110001011","111111111111101100","000000000000011001","111111111111110100","000000000000101001","000000000001101001","111111111101010101","000000000000110111","111111111101010000","111111111111111011"),
("111111111110110011","000000000000001010","000000000000000111","000000000001000100","000000000000001100","000000000001000101","000000000000010011","111111111111010111","111111111111010111","111111111111010100"),
("000000000000000110","111111111111000101","111111111111011100","000000000000011101","000000000000011100","111111111111101110","000000000001010011","111111111111011011","000000000000011011","000000000000011101"),
("111111111111010000","000000000001001111","111111111111111010","000000000001011011","000000000000000010","111111111101011011","111111111111111000","000000000000101100","111111111111001100","111111111110111001"),
("111111111111101111","000000000001101111","111111111111011000","111111111110010011","000000000001000000","000000000000000101","000000000000111101","000000000000010110","111111111110101010","111111111111001101"),
("000000000000101001","111111111110101101","111111111111011011","000000000000011011","111111111110110100","111111111111111111","000000000000001001","111111111110110101","000000000000100010","000000000000011100"),
("111111111111111101","111111111101000010","111111111111011001","111111111110010111","111111111110001000","000000000010100001","000000000001101000","000000000000001000","000000000000010000","000000000000000111"),
("000000000000111001","000000000001111000","000000000000100001","111111111111101001","000000000000000001","111111111110100010","000000000000011010","111111111110110011","111111111111100010","111111111111101111"),
("000000000000011011","111111111110101000","111111111111110010","111111111110111101","111111111111111000","111111111110110101","111111111110010101","000000000000011000","000000000000101010","000000000001000000"),
("111111111111001111","111111111101100001","111111111110000100","000000000000001110","111111111110110011","000000000000011101","111111111111101101","111111111110110101","111111111111101100","000000000001100010"),
("111111111110100101","111111111111110000","000000000000010011","000000000001111011","111111111110111111","111111111111010101","111111111110011100","111111111110110010","000000000000000101","000000000001001010"),
("111111111111100100","111111111110000111","000000000000011010","000000000000011001","000000000000000001","000000000000011000","000000000000100010","000000000000001100","000000000000010111","000000000000100011"),
("111111111111000111","000000000000010111","111111111110010010","000000000000010011","000000000000010000","000000000001100000","000000000001000100","111111111111010100","111111111110011100","111111111100111111"),
("111111111111011001","111111111111011111","111111111111010001","000000000001000110","000000000001000011","111111111101001111","111111111111101010","000000000001101110","000000000000000110","000000000000101110"),
("111111111111110100","111111111111001111","000000000001000101","111111111111010111","000000000000010101","000000000000011010","000000000000110011","111111111110010011","000000000000010011","000000000000100000"),
("111111111111100101","111111111111001100","111111111110111110","111111111110001000","000000000000100100","000000000000100110","000000000000011011","111111111110011101","000000000001100010","111111111111011001"),
("000000000000111110","111111111111001101","111111111111111101","000000000000110111","111111111110011110","000000000000000001","000000000000100111","111111111110111010","000000000000011100","000000000000110010"),
("111111111111110111","000000000000100001","000000000000001000","000000000000000100","111111111111011111","111111111111111001","111111111111100101","111111111110100001","000000000000111000","111111111111011100"),
("111111111111101101","000000000000101010","111111111111111110","111111111110010110","111111111111110001","000000000000011000","111111111111011111","000000000000100011","000000000000110111","111111111110111100"),
("000000000000101101","000000000000000010","000000000000110011","000000000000000000","111111111111101011","111111111111010100","000000000000001000","111111111111000101","000000000000111100","111111111111000110"),
("111111111111011111","111111111111111101","111111111111000101","111111111111110000","000000000000011100","111111111111010100","111111111110010111","000000000000000100","000000000000011110","000000000000111111"),
("111111111111100101","111111111110100000","111111111111101100","111111111111111000","111111111111011110","111111111101111011","000000000001100010","000000000000100111","000000000000101011","000000000000010011"),
("111111111111101000","000000000000110100","111111111110010101","000000000001000000","000000000001000111","111111111110110111","111111111110110000","000000000000000000","111111111110101110","000000000000111101"),
("000000000000110011","111111111111000000","000000000000010001","111111111110111111","000000000000100011","111111111111110011","000000000000001100","000000000000011100","111111111111110001","000000000000010011"),
("111111111111110000","000000000000000000","111111111111111000","111111111111111010","000000000000001100","111111111111101110","111111111110111011","000000000000010110","000000000000101011","000000000000100011"),
("000000000001000010","000000000001001000","000000000001001100","111111111110110110","000000000000110001","000000000000011010","111111111111011101","111111111110110101","111111111101110111","000000000001010100"),
("111111111111100011","111111111111010111","111111111111110101","000000000000010001","000000000000001000","000000000000000001","000000000000111100","111111111110111011","000000000000101111","111111111111011000"),
("111111111111100001","111111111111011110","111111111111011010","000000000000110111","000000000000000111","111111111111111001","111111111111010101","000000000000001100","000000000000100111","111111111111011101"),
("111111111110011101","111111111111100001","000000000000001100","000000000001001010","000000000000100110","111111111111010101","111111111110001110","000000000000011000","000000000000101111","000000000000000000"),
("000000000001000101","111111111111101100","000000000001000010","000000000000010110","111111111110101001","111111111110100001","000000000000011011","111111111111001101","111111111111110111","000000000001001010"),
("000000000000001110","111111111111011000","000000000000010010","000000000000110000","111111111111101101","000000000000000111","000000000000110100","111111111111110100","000000000000011110","000000000000001100"),
("000000000000011100","000000000000011111","000000000000100010","000000000000101001","111111111110110001","000000000001000001","111111111110000010","000000000000010100","111111111110111100","111111111111001000"),
("111111111111110101","000000000000000101","111111111110001010","111111111111111011","000000000000111101","000000000000101101","111111111110010101","111111111111010000","000000000000000000","000000000000110111"),
("000000000000000101","111111111111111110","000000000000000101","000000000000111101","111111111110011010","000000000000100110","111111111110011101","000000000000000000","111111111111110001","000000000000000101"),
("111111111111011111","111111111111001100","000000000000011101","111111111111101010","111111111110101000","000000000001000100","000000000000010100","000000000000100011","111111111111000110","111111111110001101"),
("000000000000011111","000000000000011000","000000000000101000","111111111110100011","000000000000100111","000000000000101011","000000000000010101","111111111111110000","000000000000001100","111111111111110011"),
("111111111111101001","000000000000000101","000000000001001000","111111111110000011","111111111111101000","111111111110111111","000000000000010010","000000000000011001","111111111111011011","000000000000100101"),
("111111111101110100","000000000010000101","000000000010100111","111111111111000010","111111111111110011","111111111110100101","000000000000101011","000000000001101111","000000000000100111","111111111101101101"),
("000000000000111100","000000000000001001","000000000001011100","111111111111100111","000000000000100111","111111111111110111","000000000000111011","000000000000101100","111111111101110111","111111111111010100"),
("000000000000101111","111111111111110010","111111111111101011","111111111111011000","111111111110001110","000000000000101100","000000000001010010","111111111111001110","000000000000000110","000000000000101000"),
("000000000000000000","111111111111000000","000000000000101100","111111111111010001","111111111101111011","000000000000001110","000000000000011000","000000000000101101","111111111111111000","111111111110111011"),
("111111111111011101","000000000000001010","111111111111001010","000000000000100000","000000000000100100","000000000000000110","111111111110101101","000000000000000000","111111111111111010","000000000000111110"));
  

constant bias_1 : intermediate_output := ("000000000000100010","111111111111101000","000000000000101011","111111111111110010","000000000000010010","000000000000011100","111111111111111111","000000000000000110","111111111111111010","000000000000000111","000000000000001100","111111111111111010","000000000000001100","000000000000011100","000000000000011100","000000000000010110","111111111111111111","000000000000001000","111111111111111100","000000000000000101","000000000000100000","000000000000001100","111111111111111110","111111111111111101","000000000000010001","000000000000001011","000000000000100010","111111111111110011","000000000000000011","000000000000001011","000000000000100000","111111111111111110","111111111111110110","111111111111111101","000000000000011101","111111111111111100","000000000000011100","000000000000010011","000000000000010001","000000000000010000","000000000000010011","000000000000011101","000000000000001100","000000000000000100","000000000000001010","000000000000000101","111111111111101001","000000000000100001","000000000000001100","111111111111100100","111111111111110100","000000000000001010","000000000000000010","000000000000000100","000000000000000111","000000000000100000","000000000000001010","111111111111101001","111111111111101110","111111111111111101","111111111111101110","000000000000001101","111111111111111011","111111111111110001","000000000000010001","000000000000010010","000000000000010111","111111111111101101","000000000000000001","000000000000100000","111111111111110100","111111111111111001","000000000000001010","111111111111111001","000000000000000000","000000000000001011","000000000000100010","111111111111101101","000000000000001011","111111111111110111","000000000000000110","111111111111110111","000000000000011010","000000000000001101","111111111111111011","000000000000000110","000000000000100000","000000000000010010","111111111111110100","111111111111111010","000000000000010011","111111111111010110","000000000000001100","111111111111111010","111111111111111111","000000000000000001","000000000000000001","000000000000001010","111111111111111101","111111111111111010","000000000000010001","000000000000000100","111111111111011110","111111111111111010","000000000000010011","111111111111110101","000000000000000000","000000000000000001","000000000000000000","000000000000011001","111111111111111111","000000000000001000","111111111111111111","111111111111110011","000000000000001011","111111111111100011","111111111111100010","000000000000000111","000000000000001111","111111111111111000","000000000000010011","000000000000100111","000000000000010100","000000000000010101","000000000000001011","111111111111110001","000000000000010101","000000000000000111");
constant bias_2 : final_output := ("111111111111011110","000000000000000110","000000000000010011","111111111111101001","000000000000001101","000000000000011110","111111111111110011","000000000000000111","111111111111111100","111111111111110101");

end package;